// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition"

// DATE "09/26/2021 10:09:45"

// 
// Device: Altera 10M50DAF484C7G Package FBGA484
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module ADC (
	altera_reserved_tms,
	altera_reserved_tck,
	altera_reserved_tdi,
	altera_reserved_tdo,
	clk_clk,
	reset_reset_n)/* synthesis synthesis_greybox=1 */;
input 	altera_reserved_tms;
input 	altera_reserved_tck;
input 	altera_reserved_tdi;
output 	altera_reserved_tdo;
input 	clk_clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \pll|sd1|wire_pll7_locked ;
wire \pll|sd1|wire_pll7_clk[0] ;
wire \avalonbridge|jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|jtag_streaming|tdo~1_combout ;
wire \adc|sample_store_internal|readdata[0]~q ;
wire \adc|sequencer_internal|u_seq_csr|readdata[0]~q ;
wire \mm_interconnect_0|adc_sample_store_csr_translator|read_latency_shift_reg[1]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[0]~combout ;
wire \mm_interconnect_0|adc_sequencer_csr_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|adc_sample_store_csr_agent_rsp_fifo|mem_used[2]~q ;
wire \avalonbridge|transacto|p2m|address[7]~q ;
wire \avalonbridge|transacto|p2m|address[6]~q ;
wire \avalonbridge|transacto|p2m|address[5]~q ;
wire \avalonbridge|transacto|p2m|address[4]~q ;
wire \mm_interconnect_0|router|Equal0~0_combout ;
wire \avalonbridge|transacto|p2m|address[9]~q ;
wire \avalonbridge|transacto|p2m|address[3]~q ;
wire \avalonbridge|transacto|p2m|address[8]~q ;
wire \mm_interconnect_0|avalonbridge_master_agent|hold_waitrequest~q ;
wire \avalonbridge|transacto|p2m|write~q ;
wire \mm_interconnect_0|avalonbridge_master_agent|av_waitrequest~1_combout ;
wire \adc|sequencer_internal|u_seq_csr|readdata[2]~q ;
wire \adc|sample_store_internal|readdata[2]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[2]~combout ;
wire \adc|sequencer_internal|u_seq_csr|readdata[1]~q ;
wire \adc|sample_store_internal|readdata[1]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[1]~combout ;
wire \adc|sample_store_internal|readdata[5]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~0_combout ;
wire \adc|sample_store_internal|readdata[7]~q ;
wire \adc|sample_store_internal|readdata[6]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~1_combout ;
wire \adc|sample_store_internal|readdata[4]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~2_combout ;
wire \adc|sequencer_internal|u_seq_csr|readdata[3]~q ;
wire \adc|sample_store_internal|readdata[3]~q ;
wire \mm_interconnect_0|rsp_mux|src_data[3]~combout ;
wire \adc|sample_store_internal|readdata[8]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~3_combout ;
wire \rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \avalonbridge|transacto|p2m|read~q ;
wire \mm_interconnect_0|cmd_demux|src1_valid~0_combout ;
wire \avalonbridge|transacto|p2m|address[2]~q ;
wire \mm_interconnect_0|rsp_mux|WideOr1~combout ;
wire \mm_interconnect_0|adc_sample_store_csr_agent_rsp_fifo|write~1_combout ;
wire \adc|sample_store_internal|readdata[10]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~4_combout ;
wire \adc|sample_store_internal|readdata[9]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~5_combout ;
wire \adc|sample_store_internal|readdata[13]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~6_combout ;
wire \adc|sample_store_internal|readdata[15]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~7_combout ;
wire \adc|sample_store_internal|readdata[14]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~8_combout ;
wire \adc|sample_store_internal|readdata[12]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~9_combout ;
wire \adc|sample_store_internal|readdata[11]~q ;
wire \mm_interconnect_0|rsp_mux|src_payload~10_combout ;
wire \avalonbridge|transacto|p2m|writedata[0]~q ;
wire \avalonbridge|transacto|p2m|writedata[2]~q ;
wire \avalonbridge|transacto|p2m|writedata[1]~q ;
wire \avalonbridge|transacto|p2m|writedata[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ;
wire \auto_hub|~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ;
wire \clk_clk~input_o ;
wire \reset_reset_n~input_o ;
wire \altera_reserved_tms~input_o ;
wire \altera_reserved_tck~input_o ;
wire \altera_reserved_tdi~input_o ;
wire \altera_internal_jtag~TCKUTAP ;
wire \altera_internal_jtag~TMSUTAP ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ;
wire \altera_internal_jtag~TDIUTAP ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ;
wire \~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~7_combout ;
wire \~QIC_CREATED_GND~I_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~15_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~14_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~23_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~17 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~15_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~19 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~22_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~12 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~14_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~12 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~14 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~6 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~8 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~21_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~22_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~19_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~20_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ;
wire \altera_internal_jtag~TDO ;


ADC_ADC_PLL pll(
	.wire_pll7_locked(\pll|sd1|wire_pll7_locked ),
	.wire_pll7_clk_0(\pll|sd1|wire_pll7_clk[0] ),
	.clk_clk(\clk_clk~input_o ));

ADC_ADC_mm_interconnect_0 mm_interconnect_0(
	.readdata_0(\adc|sample_store_internal|readdata[0]~q ),
	.readdata_01(\adc|sequencer_internal|u_seq_csr|readdata[0]~q ),
	.read_latency_shift_reg_1(\mm_interconnect_0|adc_sample_store_csr_translator|read_latency_shift_reg[1]~q ),
	.src_data_0(\mm_interconnect_0|rsp_mux|src_data[0]~combout ),
	.mem_used_1(\mm_interconnect_0|adc_sequencer_csr_agent_rsp_fifo|mem_used[1]~q ),
	.mem_used_2(\mm_interconnect_0|adc_sample_store_csr_agent_rsp_fifo|mem_used[2]~q ),
	.address_7(\avalonbridge|transacto|p2m|address[7]~q ),
	.address_6(\avalonbridge|transacto|p2m|address[6]~q ),
	.address_5(\avalonbridge|transacto|p2m|address[5]~q ),
	.address_4(\avalonbridge|transacto|p2m|address[4]~q ),
	.Equal0(\mm_interconnect_0|router|Equal0~0_combout ),
	.address_9(\avalonbridge|transacto|p2m|address[9]~q ),
	.address_3(\avalonbridge|transacto|p2m|address[3]~q ),
	.address_8(\avalonbridge|transacto|p2m|address[8]~q ),
	.hold_waitrequest(\mm_interconnect_0|avalonbridge_master_agent|hold_waitrequest~q ),
	.write(\avalonbridge|transacto|p2m|write~q ),
	.av_waitrequest(\mm_interconnect_0|avalonbridge_master_agent|av_waitrequest~1_combout ),
	.readdata_2(\adc|sequencer_internal|u_seq_csr|readdata[2]~q ),
	.readdata_21(\adc|sample_store_internal|readdata[2]~q ),
	.src_data_2(\mm_interconnect_0|rsp_mux|src_data[2]~combout ),
	.readdata_1(\adc|sequencer_internal|u_seq_csr|readdata[1]~q ),
	.readdata_11(\adc|sample_store_internal|readdata[1]~q ),
	.src_data_1(\mm_interconnect_0|rsp_mux|src_data[1]~combout ),
	.readdata_5(\adc|sample_store_internal|readdata[5]~q ),
	.src_payload(\mm_interconnect_0|rsp_mux|src_payload~0_combout ),
	.readdata_6(\adc|sample_store_internal|readdata[6]~q ),
	.src_payload1(\mm_interconnect_0|rsp_mux|src_payload~1_combout ),
	.readdata_4(\adc|sample_store_internal|readdata[4]~q ),
	.src_payload2(\mm_interconnect_0|rsp_mux|src_payload~2_combout ),
	.readdata_3(\adc|sequencer_internal|u_seq_csr|readdata[3]~q ),
	.readdata_31(\adc|sample_store_internal|readdata[3]~q ),
	.src_data_3(\mm_interconnect_0|rsp_mux|src_data[3]~combout ),
	.readdata_8(\adc|sample_store_internal|readdata[8]~q ),
	.src_payload3(\mm_interconnect_0|rsp_mux|src_payload~3_combout ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.read(\avalonbridge|transacto|p2m|read~q ),
	.src1_valid(\mm_interconnect_0|cmd_demux|src1_valid~0_combout ),
	.WideOr1(\mm_interconnect_0|rsp_mux|WideOr1~combout ),
	.write1(\mm_interconnect_0|adc_sample_store_csr_agent_rsp_fifo|write~1_combout ),
	.readdata_10(\adc|sample_store_internal|readdata[10]~q ),
	.src_payload4(\mm_interconnect_0|rsp_mux|src_payload~4_combout ),
	.readdata_9(\adc|sample_store_internal|readdata[9]~q ),
	.src_payload5(\mm_interconnect_0|rsp_mux|src_payload~5_combout ),
	.readdata_13(\adc|sample_store_internal|readdata[13]~q ),
	.src_payload6(\mm_interconnect_0|rsp_mux|src_payload~6_combout ),
	.readdata_15(\adc|sample_store_internal|readdata[15]~q ),
	.src_payload7(\mm_interconnect_0|rsp_mux|src_payload~7_combout ),
	.readdata_14(\adc|sample_store_internal|readdata[14]~q ),
	.src_payload8(\mm_interconnect_0|rsp_mux|src_payload~8_combout ),
	.readdata_12(\adc|sample_store_internal|readdata[12]~q ),
	.src_payload9(\mm_interconnect_0|rsp_mux|src_payload~9_combout ),
	.readdata_111(\adc|sample_store_internal|readdata[11]~q ),
	.src_payload10(\mm_interconnect_0|rsp_mux|src_payload~10_combout ),
	.clk_clk(\clk_clk~input_o ));

ADC_altera_reset_controller_1 rst_controller(
	.altera_reset_synchronizer_int_chain_out(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.clk_clk(\clk_clk~input_o ),
	.reset_reset_n(\reset_reset_n~input_o ));

ADC_ADC_AvalonBridge avalonbridge(
	.tdo(\avalonbridge|jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|jtag_streaming|tdo~1_combout ),
	.read_latency_shift_reg_1(\mm_interconnect_0|adc_sample_store_csr_translator|read_latency_shift_reg[1]~q ),
	.src_data_0(\mm_interconnect_0|rsp_mux|src_data[0]~combout ),
	.address_7(\avalonbridge|transacto|p2m|address[7]~q ),
	.address_6(\avalonbridge|transacto|p2m|address[6]~q ),
	.address_5(\avalonbridge|transacto|p2m|address[5]~q ),
	.address_4(\avalonbridge|transacto|p2m|address[4]~q ),
	.address_9(\avalonbridge|transacto|p2m|address[9]~q ),
	.address_3(\avalonbridge|transacto|p2m|address[3]~q ),
	.address_8(\avalonbridge|transacto|p2m|address[8]~q ),
	.master_write(\avalonbridge|transacto|p2m|write~q ),
	.av_waitrequest(\mm_interconnect_0|avalonbridge_master_agent|av_waitrequest~1_combout ),
	.src_data_2(\mm_interconnect_0|rsp_mux|src_data[2]~combout ),
	.src_data_1(\mm_interconnect_0|rsp_mux|src_data[1]~combout ),
	.src_payload(\mm_interconnect_0|rsp_mux|src_payload~0_combout ),
	.readdata_7(\adc|sample_store_internal|readdata[7]~q ),
	.src_payload1(\mm_interconnect_0|rsp_mux|src_payload~1_combout ),
	.src_payload2(\mm_interconnect_0|rsp_mux|src_payload~2_combout ),
	.src_data_3(\mm_interconnect_0|rsp_mux|src_data[3]~combout ),
	.src_payload3(\mm_interconnect_0|rsp_mux|src_payload~3_combout ),
	.master_read(\avalonbridge|transacto|p2m|read~q ),
	.address_2(\avalonbridge|transacto|p2m|address[2]~q ),
	.WideOr1(\mm_interconnect_0|rsp_mux|WideOr1~combout ),
	.src_payload4(\mm_interconnect_0|rsp_mux|src_payload~4_combout ),
	.src_payload5(\mm_interconnect_0|rsp_mux|src_payload~5_combout ),
	.src_payload6(\mm_interconnect_0|rsp_mux|src_payload~6_combout ),
	.src_payload7(\mm_interconnect_0|rsp_mux|src_payload~7_combout ),
	.src_payload8(\mm_interconnect_0|rsp_mux|src_payload~8_combout ),
	.src_payload9(\mm_interconnect_0|rsp_mux|src_payload~9_combout ),
	.src_payload10(\mm_interconnect_0|rsp_mux|src_payload~10_combout ),
	.writedata_0(\avalonbridge|transacto|p2m|writedata[0]~q ),
	.writedata_2(\avalonbridge|transacto|p2m|writedata[2]~q ),
	.writedata_1(\avalonbridge|transacto|p2m|writedata[1]~q ),
	.writedata_3(\avalonbridge|transacto|p2m|writedata[3]~q ),
	.altera_internal_jtag(\altera_internal_jtag~TCKUTAP ),
	.altera_internal_jtag1(\altera_internal_jtag~TDIUTAP ),
	.state_4(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.splitter_nodes_receive_0_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.virtual_ir_scan_reg(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.state_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.state_8(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.irf_reg_0_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.irf_reg_1_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.irf_reg_2_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][2]~q ),
	.clk_clk(\clk_clk~input_o ),
	.reset_reset_n(\reset_reset_n~input_o ));

ADC_ADC_ADC adc(
	.wire_pll7_locked(\pll|sd1|wire_pll7_locked ),
	.wire_pll7_clk_0(\pll|sd1|wire_pll7_clk[0] ),
	.readdata_0(\adc|sample_store_internal|readdata[0]~q ),
	.readdata_01(\adc|sequencer_internal|u_seq_csr|readdata[0]~q ),
	.mem_used_1(\mm_interconnect_0|adc_sequencer_csr_agent_rsp_fifo|mem_used[1]~q ),
	.mem_used_2(\mm_interconnect_0|adc_sample_store_csr_agent_rsp_fifo|mem_used[2]~q ),
	.address_7(\avalonbridge|transacto|p2m|address[7]~q ),
	.address_6(\avalonbridge|transacto|p2m|address[6]~q ),
	.address_5(\avalonbridge|transacto|p2m|address[5]~q ),
	.address_4(\avalonbridge|transacto|p2m|address[4]~q ),
	.Equal0(\mm_interconnect_0|router|Equal0~0_combout ),
	.address_3(\avalonbridge|transacto|p2m|address[3]~q ),
	.address_8(\avalonbridge|transacto|p2m|address[8]~q ),
	.hold_waitrequest(\mm_interconnect_0|avalonbridge_master_agent|hold_waitrequest~q ),
	.write(\avalonbridge|transacto|p2m|write~q ),
	.readdata_2(\adc|sequencer_internal|u_seq_csr|readdata[2]~q ),
	.readdata_21(\adc|sample_store_internal|readdata[2]~q ),
	.readdata_1(\adc|sequencer_internal|u_seq_csr|readdata[1]~q ),
	.readdata_11(\adc|sample_store_internal|readdata[1]~q ),
	.readdata_5(\adc|sample_store_internal|readdata[5]~q ),
	.readdata_7(\adc|sample_store_internal|readdata[7]~q ),
	.readdata_6(\adc|sample_store_internal|readdata[6]~q ),
	.readdata_4(\adc|sample_store_internal|readdata[4]~q ),
	.readdata_3(\adc|sequencer_internal|u_seq_csr|readdata[3]~q ),
	.readdata_31(\adc|sample_store_internal|readdata[3]~q ),
	.readdata_8(\adc|sample_store_internal|readdata[8]~q ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.read(\avalonbridge|transacto|p2m|read~q ),
	.src1_valid(\mm_interconnect_0|cmd_demux|src1_valid~0_combout ),
	.address_2(\avalonbridge|transacto|p2m|address[2]~q ),
	.write1(\mm_interconnect_0|adc_sample_store_csr_agent_rsp_fifo|write~1_combout ),
	.readdata_10(\adc|sample_store_internal|readdata[10]~q ),
	.readdata_9(\adc|sample_store_internal|readdata[9]~q ),
	.readdata_13(\adc|sample_store_internal|readdata[13]~q ),
	.readdata_15(\adc|sample_store_internal|readdata[15]~q ),
	.readdata_14(\adc|sample_store_internal|readdata[14]~q ),
	.readdata_12(\adc|sample_store_internal|readdata[12]~q ),
	.readdata_111(\adc|sample_store_internal|readdata[11]~q ),
	.writedata_0(\avalonbridge|transacto|p2m|writedata[0]~q ),
	.writedata_2(\avalonbridge|transacto|p2m|writedata[2]~q ),
	.writedata_1(\avalonbridge|transacto|p2m|writedata[1]~q ),
	.writedata_3(\avalonbridge|transacto|p2m|writedata[3]~q ),
	.GND_port(\~GND~combout ),
	.clk_clk(\clk_clk~input_o ));

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][2] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .lut_mask = 16'hEFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .lut_mask = 16'hFAFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .lut_mask = 16'hB8FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .sum_lutc_input = "datac";

assign \clk_clk~input_o  = clk_clk;

assign \reset_reset_n~input_o  = reset_reset_n;

assign altera_reserved_tdo = \altera_internal_jtag~TDO ;

assign \altera_reserved_tms~input_o  = altera_reserved_tms;

assign \altera_reserved_tck~input_o  = altera_reserved_tck;

assign \altera_reserved_tdi~input_o  = altera_reserved_tdi;

fiftyfivenm_jtag altera_internal_jtag(
	.tms(\altera_reserved_tms~input_o ),
	.tck(\altera_reserved_tck~input_o ),
	.tdi(\altera_reserved_tdi~input_o ),
	.tdouser(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.tdo(\altera_internal_jtag~TDO ),
	.tmsutap(\altera_internal_jtag~TMSUTAP ),
	.tckutap(\altera_internal_jtag~TCKUTAP ),
	.tdiutap(\altera_internal_jtag~TDIUTAP ),
	.shiftuser(),
	.clkdruser(),
	.updateuser(),
	.runidleuser(),
	.usr1user());

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\altera_internal_jtag~TMSUTAP ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .lut_mask = 16'h0FF0;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .lut_mask = 16'hC33C;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .lut_mask = 16'hFF7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\altera_internal_jtag~TMSUTAP ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\~GND~combout ),
	.cout());
defparam \~GND .lut_mask = 16'h0000;
defparam \~GND .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .lut_mask = 16'h7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~10 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~10 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~10 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~11 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~11 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~7 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~7 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \~QIC_CREATED_GND~I (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\~QIC_CREATED_GND~I_combout ),
	.cout());
defparam \~QIC_CREATED_GND~I .lut_mask = 16'h0000;
defparam \~QIC_CREATED_GND~I .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~12 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~10_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~11_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~7_combout ),
	.datad(\~QIC_CREATED_GND~I_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~12 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~12 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9 (
	.dataa(\~GND~combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~6 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~6 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~6 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~6 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~15 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~6_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~15_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~15 .lut_mask = 16'hFFAC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~15 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~9_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~15_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~8 (
	.dataa(\~GND~combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~8 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~8 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~8_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~15_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~0 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1 .lut_mask = 16'hFDFD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~2 .lut_mask = 16'h6996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~2_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3 .lut_mask = 16'hEBBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~4 .lut_mask = 16'h0FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~4 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~4_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5 .lut_mask = 16'hFAFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~5_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~12_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~5 .lut_mask = 16'hEEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~5_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~7_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~13 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~14 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~13_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~14_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~14 .lut_mask = 16'hACFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~14 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~14_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 (
	.dataa(\~GND~combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~15_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .lut_mask = 16'h3FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~12 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11 .lut_mask = 16'h55AA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~12 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~17 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16 .lut_mask = 16'h5AAF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~23 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~23_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~23 .lut_mask = 16'hFFFB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~23 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~17 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~19 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~15 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~15_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~15 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~15 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~19 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20 .lut_mask = 16'h5A5A;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~22 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~15_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~22_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~22 .lut_mask = 16'hFFEF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~22 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~14 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~14_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~14 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~14 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~14_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .lut_mask = 16'hBF8F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9 .lut_mask = 16'hAFCF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10 .lut_mask = 16'hFFEF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~14_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .lut_mask = 16'hFFF6;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .lut_mask = 16'hBF8F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~14_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~14_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .lut_mask = 16'hD8FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~6 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5 .lut_mask = 16'h55AA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~8 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~11_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~12 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~11 .lut_mask = 16'h5AAF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~11 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~12 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~14 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~10 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~10 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~9_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~10_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~14 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15 .lut_mask = 16'h5A5A;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~9_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~10_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 .lut_mask = 16'h0FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13 .lut_mask = 16'h0FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~9 .lut_mask = 16'hFFFD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~9 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~9_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~10_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~6 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~7_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~8 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~7 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~7 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~9_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~10_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~9_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~10_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~21 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~21_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~21 .lut_mask = 16'h6996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~21 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~22 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~21_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~22_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~22 .lut_mask = 16'hDFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~22 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1 .lut_mask = 16'hEEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~11 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~11 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~12 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~11_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~12 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~12 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~22_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~12_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~19 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~19_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~19 .lut_mask = 16'h6996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~19 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~20 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~19_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~20_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~20 .lut_mask = 16'hEDDE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~20 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~20_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~12_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14 .lut_mask = 16'hEBBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15 (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15 .lut_mask = 16'hC33C;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~16_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~12_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17 .lut_mask = 16'h7FF7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~17_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18 .lut_mask = 16'hEDDE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~18_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~12_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .lut_mask = 16'h0FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena .lut_mask = 16'hFFFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3_combout ),
	.asdata(\altera_internal_jtag~TDIUTAP ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0] .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~12 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7_combout ),
	.datad(\avalonbridge|jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|jtag_streaming|tdo~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~12 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~12 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9 .lut_mask = 16'hF7F7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~9_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10 .lut_mask = 16'hFFEF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~8_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~12_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~10_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~11 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~11 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo (
	.clk(!\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .power_up = "low";

fiftyfivenm_lcell_comb \auto_hub|~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|~GND~combout ),
	.cout());
defparam \auto_hub|~GND .lut_mask = 16'h0000;
defparam \auto_hub|~GND .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .sum_lutc_input = "datac";

endmodule

module ADC_ADC_ADC (
	wire_pll7_locked,
	wire_pll7_clk_0,
	readdata_0,
	readdata_01,
	mem_used_1,
	mem_used_2,
	address_7,
	address_6,
	address_5,
	address_4,
	Equal0,
	address_3,
	address_8,
	hold_waitrequest,
	write,
	readdata_2,
	readdata_21,
	readdata_1,
	readdata_11,
	readdata_5,
	readdata_7,
	readdata_6,
	readdata_4,
	readdata_3,
	readdata_31,
	readdata_8,
	altera_reset_synchronizer_int_chain_out,
	read,
	src1_valid,
	address_2,
	write1,
	readdata_10,
	readdata_9,
	readdata_13,
	readdata_15,
	readdata_14,
	readdata_12,
	readdata_111,
	writedata_0,
	writedata_2,
	writedata_1,
	writedata_3,
	GND_port,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_locked;
input 	wire_pll7_clk_0;
output 	readdata_0;
output 	readdata_01;
input 	mem_used_1;
input 	mem_used_2;
input 	address_7;
input 	address_6;
input 	address_5;
input 	address_4;
input 	Equal0;
input 	address_3;
input 	address_8;
input 	hold_waitrequest;
input 	write;
output 	readdata_2;
output 	readdata_21;
output 	readdata_1;
output 	readdata_11;
output 	readdata_5;
output 	readdata_7;
output 	readdata_6;
output 	readdata_4;
output 	readdata_3;
output 	readdata_31;
output 	readdata_8;
input 	altera_reset_synchronizer_int_chain_out;
input 	read;
input 	src1_valid;
input 	address_2;
input 	write1;
output 	readdata_10;
output 	readdata_9;
output 	readdata_13;
output 	readdata_15;
output 	readdata_14;
output 	readdata_12;
output 	readdata_111;
input 	writedata_0;
input 	writedata_2;
input 	writedata_1;
input 	writedata_3;
input 	GND_port;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \control_internal|u_control_fsm|rsp_valid~q ;
wire \control_internal|u_control_fsm|rsp_data[0]~q ;
wire \control_internal|u_control_fsm|cmd_ready~q ;
wire \control_internal|u_control_fsm|rsp_data[2]~q ;
wire \control_internal|u_control_fsm|rsp_data[1]~q ;
wire \control_internal|u_control_fsm|rsp_data[5]~q ;
wire \control_internal|u_control_fsm|rsp_data[7]~q ;
wire \control_internal|u_control_fsm|rsp_data[6]~q ;
wire \control_internal|u_control_fsm|rsp_data[4]~q ;
wire \control_internal|u_control_fsm|rsp_data[3]~q ;
wire \control_internal|u_control_fsm|rsp_data[8]~q ;
wire \sequencer_internal|u_seq_ctrl|cmd_channel[4]~q ;
wire \control_internal|u_control_fsm|rsp_eop~q ;
wire \control_internal|u_control_fsm|rsp_data[10]~q ;
wire \control_internal|u_control_fsm|rsp_data[9]~q ;
wire \control_internal|u_control_fsm|rsp_data[11]~q ;
wire \sequencer_internal|u_seq_ctrl|cmd_eop~q ;


ADC_altera_modular_adc_sequencer sequencer_internal(
	.readdata_0(readdata_01),
	.mem_used_1(mem_used_1),
	.write(write),
	.readdata_2(readdata_2),
	.readdata_1(readdata_1),
	.readdata_3(readdata_3),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.read(read),
	.src1_valid(src1_valid),
	.address_2(address_2),
	.cmd_ready(\control_internal|u_control_fsm|cmd_ready~q ),
	.writedata_0(writedata_0),
	.writedata_2(writedata_2),
	.writedata_1(writedata_1),
	.writedata_3(writedata_3),
	.cmd_channel_4(\sequencer_internal|u_seq_ctrl|cmd_channel[4]~q ),
	.cmd_eop(\sequencer_internal|u_seq_ctrl|cmd_eop~q ),
	.clk_clk(clk_clk));

ADC_altera_modular_adc_sample_store sample_store_internal(
	.readdata_0(readdata_0),
	.mem_used_2(mem_used_2),
	.address_7(address_7),
	.address_6(address_6),
	.address_5(address_5),
	.address_4(address_4),
	.Equal0(Equal0),
	.address_3(address_3),
	.address_8(address_8),
	.hold_waitrequest(hold_waitrequest),
	.write(write),
	.readdata_2(readdata_21),
	.readdata_1(readdata_11),
	.readdata_5(readdata_5),
	.readdata_7(readdata_7),
	.readdata_6(readdata_6),
	.readdata_4(readdata_4),
	.readdata_3(readdata_31),
	.readdata_8(readdata_8),
	.rst_n(altera_reset_synchronizer_int_chain_out),
	.address_2(address_2),
	.write1(write1),
	.readdata_10(readdata_10),
	.readdata_9(readdata_9),
	.readdata_13(readdata_13),
	.readdata_15(readdata_15),
	.readdata_14(readdata_14),
	.readdata_12(readdata_12),
	.readdata_11(readdata_111),
	.rsp_valid(\control_internal|u_control_fsm|rsp_valid~q ),
	.rsp_data_0(\control_internal|u_control_fsm|rsp_data[0]~q ),
	.writedata_0(writedata_0),
	.rsp_data_2(\control_internal|u_control_fsm|rsp_data[2]~q ),
	.rsp_data_1(\control_internal|u_control_fsm|rsp_data[1]~q ),
	.rsp_data_5(\control_internal|u_control_fsm|rsp_data[5]~q ),
	.rsp_data_7(\control_internal|u_control_fsm|rsp_data[7]~q ),
	.rsp_data_6(\control_internal|u_control_fsm|rsp_data[6]~q ),
	.rsp_data_4(\control_internal|u_control_fsm|rsp_data[4]~q ),
	.rsp_data_3(\control_internal|u_control_fsm|rsp_data[3]~q ),
	.rsp_data_8(\control_internal|u_control_fsm|rsp_data[8]~q ),
	.rsp_eop(\control_internal|u_control_fsm|rsp_eop~q ),
	.rsp_data_10(\control_internal|u_control_fsm|rsp_data[10]~q ),
	.rsp_data_9(\control_internal|u_control_fsm|rsp_data[9]~q ),
	.rsp_data_11(\control_internal|u_control_fsm|rsp_data[11]~q ),
	.GND_port(GND_port),
	.clk_clk(clk_clk));

ADC_altera_modular_adc_control control_internal(
	.wire_pll7_locked(wire_pll7_locked),
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.rsp_valid(\control_internal|u_control_fsm|rsp_valid~q ),
	.rsp_data_0(\control_internal|u_control_fsm|rsp_data[0]~q ),
	.cmd_ready(\control_internal|u_control_fsm|cmd_ready~q ),
	.rsp_data_2(\control_internal|u_control_fsm|rsp_data[2]~q ),
	.rsp_data_1(\control_internal|u_control_fsm|rsp_data[1]~q ),
	.rsp_data_5(\control_internal|u_control_fsm|rsp_data[5]~q ),
	.rsp_data_7(\control_internal|u_control_fsm|rsp_data[7]~q ),
	.rsp_data_6(\control_internal|u_control_fsm|rsp_data[6]~q ),
	.rsp_data_4(\control_internal|u_control_fsm|rsp_data[4]~q ),
	.rsp_data_3(\control_internal|u_control_fsm|rsp_data[3]~q ),
	.rsp_data_8(\control_internal|u_control_fsm|rsp_data[8]~q ),
	.cmd_channel_4(\sequencer_internal|u_seq_ctrl|cmd_channel[4]~q ),
	.rsp_eop(\control_internal|u_control_fsm|rsp_eop~q ),
	.rsp_data_10(\control_internal|u_control_fsm|rsp_data[10]~q ),
	.rsp_data_9(\control_internal|u_control_fsm|rsp_data[9]~q ),
	.rsp_data_11(\control_internal|u_control_fsm|rsp_data[11]~q ),
	.cmd_eop(\sequencer_internal|u_seq_ctrl|cmd_eop~q ),
	.GND_port(GND_port),
	.clk_clk(clk_clk));

endmodule

module ADC_altera_modular_adc_control (
	wire_pll7_locked,
	wire_pll7_clk_0,
	altera_reset_synchronizer_int_chain_out,
	rsp_valid,
	rsp_data_0,
	cmd_ready,
	rsp_data_2,
	rsp_data_1,
	rsp_data_5,
	rsp_data_7,
	rsp_data_6,
	rsp_data_4,
	rsp_data_3,
	rsp_data_8,
	cmd_channel_4,
	rsp_eop,
	rsp_data_10,
	rsp_data_9,
	rsp_data_11,
	cmd_eop,
	GND_port,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	wire_pll7_locked;
input 	wire_pll7_clk_0;
input 	altera_reset_synchronizer_int_chain_out;
output 	rsp_valid;
output 	rsp_data_0;
output 	cmd_ready;
output 	rsp_data_2;
output 	rsp_data_1;
output 	rsp_data_5;
output 	rsp_data_7;
output 	rsp_data_6;
output 	rsp_data_4;
output 	rsp_data_3;
output 	rsp_data_8;
input 	cmd_channel_4;
output 	rsp_eop;
output 	rsp_data_10;
output 	rsp_data_9;
output 	rsp_data_11;
input 	cmd_eop;
input 	GND_port;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \adc_inst|adcblock_instance|eoc ;
wire \adc_inst|adcblock_instance|clkout_adccore ;
wire \adc_inst|adcblock_instance|wire_from_adc_dout[0] ;
wire \adc_inst|adcblock_instance|wire_from_adc_dout[1] ;
wire \adc_inst|adcblock_instance|wire_from_adc_dout[2] ;
wire \adc_inst|adcblock_instance|wire_from_adc_dout[3] ;
wire \adc_inst|adcblock_instance|wire_from_adc_dout[4] ;
wire \adc_inst|adcblock_instance|wire_from_adc_dout[5] ;
wire \adc_inst|adcblock_instance|wire_from_adc_dout[6] ;
wire \adc_inst|adcblock_instance|wire_from_adc_dout[7] ;
wire \adc_inst|adcblock_instance|wire_from_adc_dout[8] ;
wire \adc_inst|adcblock_instance|wire_from_adc_dout[9] ;
wire \adc_inst|adcblock_instance|wire_from_adc_dout[10] ;
wire \adc_inst|adcblock_instance|wire_from_adc_dout[11] ;
wire \u_control_fsm|soc~q ;
wire \u_control_fsm|chsel[1]~q ;
wire \u_control_fsm|chsel[0]~q ;
wire \u_control_fsm|chsel[1]~_wirecell_combout ;
wire \u_control_fsm|usr_pwd~_wirecell_combout ;


ADC_fiftyfivenm_adcblock_top_wrapper adc_inst(
	.eoc(\adc_inst|adcblock_instance|eoc ),
	.clkout_adccore(\adc_inst|adcblock_instance|clkout_adccore ),
	.wire_from_adc_dout_0(\adc_inst|adcblock_instance|wire_from_adc_dout[0] ),
	.wire_from_adc_dout_1(\adc_inst|adcblock_instance|wire_from_adc_dout[1] ),
	.wire_from_adc_dout_2(\adc_inst|adcblock_instance|wire_from_adc_dout[2] ),
	.wire_from_adc_dout_3(\adc_inst|adcblock_instance|wire_from_adc_dout[3] ),
	.wire_from_adc_dout_4(\adc_inst|adcblock_instance|wire_from_adc_dout[4] ),
	.wire_from_adc_dout_5(\adc_inst|adcblock_instance|wire_from_adc_dout[5] ),
	.wire_from_adc_dout_6(\adc_inst|adcblock_instance|wire_from_adc_dout[6] ),
	.wire_from_adc_dout_7(\adc_inst|adcblock_instance|wire_from_adc_dout[7] ),
	.wire_from_adc_dout_8(\adc_inst|adcblock_instance|wire_from_adc_dout[8] ),
	.wire_from_adc_dout_9(\adc_inst|adcblock_instance|wire_from_adc_dout[9] ),
	.wire_from_adc_dout_10(\adc_inst|adcblock_instance|wire_from_adc_dout[10] ),
	.wire_from_adc_dout_11(\adc_inst|adcblock_instance|wire_from_adc_dout[11] ),
	.wire_pll7_clk_0(wire_pll7_clk_0),
	.soc(\u_control_fsm|soc~q ),
	.chsel_1(\u_control_fsm|chsel[1]~q ),
	.chsel_0(\u_control_fsm|chsel[0]~q ),
	.GND_port(GND_port),
	.chsel_11(\u_control_fsm|chsel[1]~_wirecell_combout ),
	.usr_pwd(\u_control_fsm|usr_pwd~_wirecell_combout ));

ADC_altera_modular_adc_control_fsm u_control_fsm(
	.eoc(\adc_inst|adcblock_instance|eoc ),
	.clkout_adccore(\adc_inst|adcblock_instance|clkout_adccore ),
	.wire_from_adc_dout_0(\adc_inst|adcblock_instance|wire_from_adc_dout[0] ),
	.wire_from_adc_dout_1(\adc_inst|adcblock_instance|wire_from_adc_dout[1] ),
	.wire_from_adc_dout_2(\adc_inst|adcblock_instance|wire_from_adc_dout[2] ),
	.wire_from_adc_dout_3(\adc_inst|adcblock_instance|wire_from_adc_dout[3] ),
	.wire_from_adc_dout_4(\adc_inst|adcblock_instance|wire_from_adc_dout[4] ),
	.wire_from_adc_dout_5(\adc_inst|adcblock_instance|wire_from_adc_dout[5] ),
	.wire_from_adc_dout_6(\adc_inst|adcblock_instance|wire_from_adc_dout[6] ),
	.wire_from_adc_dout_7(\adc_inst|adcblock_instance|wire_from_adc_dout[7] ),
	.wire_from_adc_dout_8(\adc_inst|adcblock_instance|wire_from_adc_dout[8] ),
	.wire_from_adc_dout_9(\adc_inst|adcblock_instance|wire_from_adc_dout[9] ),
	.wire_from_adc_dout_10(\adc_inst|adcblock_instance|wire_from_adc_dout[10] ),
	.wire_from_adc_dout_11(\adc_inst|adcblock_instance|wire_from_adc_dout[11] ),
	.wire_pll7_locked(wire_pll7_locked),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.rsp_valid1(rsp_valid),
	.rsp_data_0(rsp_data_0),
	.cmd_ready1(cmd_ready),
	.rsp_data_2(rsp_data_2),
	.rsp_data_1(rsp_data_1),
	.rsp_data_5(rsp_data_5),
	.rsp_data_7(rsp_data_7),
	.rsp_data_6(rsp_data_6),
	.rsp_data_4(rsp_data_4),
	.rsp_data_3(rsp_data_3),
	.rsp_data_8(rsp_data_8),
	.cmd_channel_4(cmd_channel_4),
	.rsp_eop1(rsp_eop),
	.rsp_data_10(rsp_data_10),
	.rsp_data_9(rsp_data_9),
	.rsp_data_11(rsp_data_11),
	.soc1(\u_control_fsm|soc~q ),
	.chsel_1(\u_control_fsm|chsel[1]~q ),
	.chsel_0(\u_control_fsm|chsel[0]~q ),
	.cmd_eop(cmd_eop),
	.chsel_11(\u_control_fsm|chsel[1]~_wirecell_combout ),
	.usr_pwd1(\u_control_fsm|usr_pwd~_wirecell_combout ),
	.clk_clk(clk_clk));

endmodule

module ADC_altera_modular_adc_control_fsm (
	eoc,
	clkout_adccore,
	wire_from_adc_dout_0,
	wire_from_adc_dout_1,
	wire_from_adc_dout_2,
	wire_from_adc_dout_3,
	wire_from_adc_dout_4,
	wire_from_adc_dout_5,
	wire_from_adc_dout_6,
	wire_from_adc_dout_7,
	wire_from_adc_dout_8,
	wire_from_adc_dout_9,
	wire_from_adc_dout_10,
	wire_from_adc_dout_11,
	wire_pll7_locked,
	altera_reset_synchronizer_int_chain_out,
	rsp_valid1,
	rsp_data_0,
	cmd_ready1,
	rsp_data_2,
	rsp_data_1,
	rsp_data_5,
	rsp_data_7,
	rsp_data_6,
	rsp_data_4,
	rsp_data_3,
	rsp_data_8,
	cmd_channel_4,
	rsp_eop1,
	rsp_data_10,
	rsp_data_9,
	rsp_data_11,
	soc1,
	chsel_1,
	chsel_0,
	cmd_eop,
	chsel_11,
	usr_pwd1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	eoc;
input 	clkout_adccore;
input 	wire_from_adc_dout_0;
input 	wire_from_adc_dout_1;
input 	wire_from_adc_dout_2;
input 	wire_from_adc_dout_3;
input 	wire_from_adc_dout_4;
input 	wire_from_adc_dout_5;
input 	wire_from_adc_dout_6;
input 	wire_from_adc_dout_7;
input 	wire_from_adc_dout_8;
input 	wire_from_adc_dout_9;
input 	wire_from_adc_dout_10;
input 	wire_from_adc_dout_11;
input 	wire_pll7_locked;
input 	altera_reset_synchronizer_int_chain_out;
output 	rsp_valid1;
output 	rsp_data_0;
output 	cmd_ready1;
output 	rsp_data_2;
output 	rsp_data_1;
output 	rsp_data_5;
output 	rsp_data_7;
output 	rsp_data_6;
output 	rsp_data_4;
output 	rsp_data_3;
output 	rsp_data_8;
input 	cmd_channel_4;
output 	rsp_eop1;
output 	rsp_data_10;
output 	rsp_data_9;
output 	rsp_data_11;
output 	soc1;
output 	chsel_1;
output 	chsel_0;
input 	cmd_eop;
output 	chsel_11;
output 	usr_pwd1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \u_eoc_synchronizer|dreg[0]~q ;
wire \u_clk_dft_synchronizer|dreg[0]~q ;
wire \eoc_synch_dly~q ;
wire \ctrl_state.PUTRESP_DLY2~q ;
wire \ctrl_state.PUTRESP_DLY3~q ;
wire \Selector6~1_combout ;
wire \Selector6~2_combout ;
wire \ctrl_state.WAIT~q ;
wire \ctrl_state_nxt.GETCMD_W~0_combout ;
wire \ctrl_state.GETCMD_W~q ;
wire \Selector1~0_combout ;
wire \Selector1~2_combout ;
wire \ctrl_state.PWRDWN~q ;
wire \Add0~0_combout ;
wire \int_timer~7_combout ;
wire \load_int_timer~0_combout ;
wire \Add0~13 ;
wire \Add0~14_combout ;
wire \int_timer~8_combout ;
wire \int_timer[7]~q ;
wire \Selector2~0_combout ;
wire \ctrl_state.PWRDWN_TSEN~q ;
wire \int_timer[6]~0_combout ;
wire \int_timer[0]~q ;
wire \Add0~1 ;
wire \Add0~2_combout ;
wire \int_timer~6_combout ;
wire \int_timer[1]~q ;
wire \Add0~3 ;
wire \Add0~4_combout ;
wire \int_timer~5_combout ;
wire \int_timer[2]~q ;
wire \Add0~5 ;
wire \Add0~6_combout ;
wire \int_timer~4_combout ;
wire \int_timer[3]~q ;
wire \Add0~7 ;
wire \Add0~8_combout ;
wire \int_timer~3_combout ;
wire \int_timer[4]~q ;
wire \Add0~9 ;
wire \Add0~10_combout ;
wire \int_timer~2_combout ;
wire \int_timer[5]~q ;
wire \Add0~11 ;
wire \Add0~12_combout ;
wire \int_timer[6]~1_combout ;
wire \int_timer[6]~q ;
wire \Selector0~0_combout ;
wire \ctrl_state.IDLE~q ;
wire \Selector1~1_combout ;
wire \cmd_fetched~0_combout ;
wire \Selector5~0_combout ;
wire \Selector3~0_combout ;
wire \clk_dft_synch_dly~q ;
wire \Selector3~1_combout ;
wire \ctrl_state.PWRDWN_DONE~q ;
wire \Selector4~0_combout ;
wire \ctrl_state.PWRUP_CH~q ;
wire \Selector5~1_combout ;
wire \ctrl_state.PWRUP_SOC~q ;
wire \Selector6~0_combout ;
wire \cmd_fetched~1_combout ;
wire \cmd_fetched~q ;
wire \Selector7~0_combout ;
wire \Selector7~1_combout ;
wire \ctrl_state.GETCMD~q ;
wire \Selector9~0_combout ;
wire \ctrl_state_nxt~0_combout ;
wire \Selector8~0_combout ;
wire \ctrl_state.PRE_CONV~q ;
wire \Selector9~1_combout ;
wire \ctrl_state.CONV~q ;
wire \ctrl_state_nxt.CONV_DLY1~0_combout ;
wire \ctrl_state.CONV_DLY1~q ;
wire \conv_dly1_s_flp~q ;
wire \pend~0_combout ;
wire \pend~q ;
wire \Selector11~0_combout ;
wire \Selector11~1_combout ;
wire \ctrl_state.WAIT_PEND~q ;
wire \ctrl_state_nxt.WAIT_PEND_DLY1~0_combout ;
wire \ctrl_state.WAIT_PEND_DLY1~q ;
wire \ctrl_state.PUTRESP_PEND~q ;
wire \Selector10~0_combout ;
wire \ctrl_state.PUTRESP~q ;
wire \load_rsp~combout ;
wire \load_dout~2_combout ;
wire \load_dout~3_combout ;
wire \dout_flp[0]~q ;
wire \rsp_data~0_combout ;
wire \dout_flp[2]~q ;
wire \rsp_data~1_combout ;
wire \dout_flp[1]~q ;
wire \rsp_data~2_combout ;
wire \dout_flp[5]~q ;
wire \rsp_data~3_combout ;
wire \dout_flp[7]~q ;
wire \rsp_data~4_combout ;
wire \dout_flp[6]~q ;
wire \rsp_data~5_combout ;
wire \dout_flp[4]~q ;
wire \rsp_data~6_combout ;
wire \dout_flp[3]~q ;
wire \rsp_data~7_combout ;
wire \dout_flp[8]~q ;
wire \rsp_data~8_combout ;
wire \cmd_eop_dly~0_combout ;
wire \cmd_eop_dly~q ;
wire \rsp_eop~0_combout ;
wire \dout_flp[10]~q ;
wire \rsp_data~9_combout ;
wire \dout_flp[9]~q ;
wire \rsp_data~10_combout ;
wire \dout_flp[11]~q ;
wire \rsp_data~11_combout ;
wire \WideOr12~0_combout ;
wire \WideOr12~1_combout ;
wire \WideOr12~2_combout ;
wire \WideOr12~3_combout ;
wire \WideOr13~0_combout ;
wire \WideOr15~0_combout ;
wire \Selector17~0_combout ;
wire \WideOr12~4_combout ;
wire \WideOr12~combout ;
wire \Selector15~0_combout ;
wire \Selector16~0_combout ;
wire \Selector18~0_combout ;
wire \Selector18~1_combout ;
wire \usr_pwd~q ;


ADC_altera_std_synchronizer_1 u_eoc_synchronizer(
	.din(eoc),
	.reset_n(altera_reset_synchronizer_int_chain_out),
	.dreg_0(\u_eoc_synchronizer|dreg[0]~q ),
	.clk(clk_clk));

ADC_altera_std_synchronizer u_clk_dft_synchronizer(
	.din(clkout_adccore),
	.reset_n(altera_reset_synchronizer_int_chain_out),
	.dreg_0(\u_clk_dft_synchronizer|dreg[0]~q ),
	.clk(clk_clk));

dffeas rsp_valid(
	.clk(clk_clk),
	.d(\load_rsp~combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rsp_valid1),
	.prn(vcc));
defparam rsp_valid.is_wysiwyg = "true";
defparam rsp_valid.power_up = "low";

dffeas \rsp_data[0] (
	.clk(clk_clk),
	.d(\rsp_data~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rsp_data_0),
	.prn(vcc));
defparam \rsp_data[0] .is_wysiwyg = "true";
defparam \rsp_data[0] .power_up = "low";

dffeas cmd_ready(
	.clk(clk_clk),
	.d(\ctrl_state.PUTRESP~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(cmd_ready1),
	.prn(vcc));
defparam cmd_ready.is_wysiwyg = "true";
defparam cmd_ready.power_up = "low";

dffeas \rsp_data[2] (
	.clk(clk_clk),
	.d(\rsp_data~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rsp_data_2),
	.prn(vcc));
defparam \rsp_data[2] .is_wysiwyg = "true";
defparam \rsp_data[2] .power_up = "low";

dffeas \rsp_data[1] (
	.clk(clk_clk),
	.d(\rsp_data~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rsp_data_1),
	.prn(vcc));
defparam \rsp_data[1] .is_wysiwyg = "true";
defparam \rsp_data[1] .power_up = "low";

dffeas \rsp_data[5] (
	.clk(clk_clk),
	.d(\rsp_data~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rsp_data_5),
	.prn(vcc));
defparam \rsp_data[5] .is_wysiwyg = "true";
defparam \rsp_data[5] .power_up = "low";

dffeas \rsp_data[7] (
	.clk(clk_clk),
	.d(\rsp_data~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rsp_data_7),
	.prn(vcc));
defparam \rsp_data[7] .is_wysiwyg = "true";
defparam \rsp_data[7] .power_up = "low";

dffeas \rsp_data[6] (
	.clk(clk_clk),
	.d(\rsp_data~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rsp_data_6),
	.prn(vcc));
defparam \rsp_data[6] .is_wysiwyg = "true";
defparam \rsp_data[6] .power_up = "low";

dffeas \rsp_data[4] (
	.clk(clk_clk),
	.d(\rsp_data~6_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rsp_data_4),
	.prn(vcc));
defparam \rsp_data[4] .is_wysiwyg = "true";
defparam \rsp_data[4] .power_up = "low";

dffeas \rsp_data[3] (
	.clk(clk_clk),
	.d(\rsp_data~7_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rsp_data_3),
	.prn(vcc));
defparam \rsp_data[3] .is_wysiwyg = "true";
defparam \rsp_data[3] .power_up = "low";

dffeas \rsp_data[8] (
	.clk(clk_clk),
	.d(\rsp_data~8_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rsp_data_8),
	.prn(vcc));
defparam \rsp_data[8] .is_wysiwyg = "true";
defparam \rsp_data[8] .power_up = "low";

dffeas rsp_eop(
	.clk(clk_clk),
	.d(\rsp_eop~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rsp_eop1),
	.prn(vcc));
defparam rsp_eop.is_wysiwyg = "true";
defparam rsp_eop.power_up = "low";

dffeas \rsp_data[10] (
	.clk(clk_clk),
	.d(\rsp_data~9_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rsp_data_10),
	.prn(vcc));
defparam \rsp_data[10] .is_wysiwyg = "true";
defparam \rsp_data[10] .power_up = "low";

dffeas \rsp_data[9] (
	.clk(clk_clk),
	.d(\rsp_data~10_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rsp_data_9),
	.prn(vcc));
defparam \rsp_data[9] .is_wysiwyg = "true";
defparam \rsp_data[9] .power_up = "low";

dffeas \rsp_data[11] (
	.clk(clk_clk),
	.d(\rsp_data~11_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rsp_data_11),
	.prn(vcc));
defparam \rsp_data[11] .is_wysiwyg = "true";
defparam \rsp_data[11] .power_up = "low";

dffeas soc(
	.clk(clk_clk),
	.d(\Selector17~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(soc1),
	.prn(vcc));
defparam soc.is_wysiwyg = "true";
defparam soc.power_up = "low";

dffeas \chsel[1] (
	.clk(clk_clk),
	.d(\Selector15~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(chsel_1),
	.prn(vcc));
defparam \chsel[1] .is_wysiwyg = "true";
defparam \chsel[1] .power_up = "low";

dffeas \chsel[0] (
	.clk(clk_clk),
	.d(\Selector16~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(chsel_0),
	.prn(vcc));
defparam \chsel[0] .is_wysiwyg = "true";
defparam \chsel[0] .power_up = "low";

fiftyfivenm_lcell_comb \chsel[1]~_wirecell (
	.dataa(chsel_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(chsel_11),
	.cout());
defparam \chsel[1]~_wirecell .lut_mask = 16'h5555;
defparam \chsel[1]~_wirecell .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \usr_pwd~_wirecell (
	.dataa(\usr_pwd~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(usr_pwd1),
	.cout());
defparam \usr_pwd~_wirecell .lut_mask = 16'h5555;
defparam \usr_pwd~_wirecell .sum_lutc_input = "datac";

dffeas eoc_synch_dly(
	.clk(clk_clk),
	.d(\u_eoc_synchronizer|dreg[0]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\eoc_synch_dly~q ),
	.prn(vcc));
defparam eoc_synch_dly.is_wysiwyg = "true";
defparam eoc_synch_dly.power_up = "low";

dffeas \ctrl_state.PUTRESP_DLY2 (
	.clk(clk_clk),
	.d(cmd_ready1),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_state.PUTRESP_DLY2~q ),
	.prn(vcc));
defparam \ctrl_state.PUTRESP_DLY2 .is_wysiwyg = "true";
defparam \ctrl_state.PUTRESP_DLY2 .power_up = "low";

dffeas \ctrl_state.PUTRESP_DLY3 (
	.clk(clk_clk),
	.d(\ctrl_state.PUTRESP_DLY2~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_state.PUTRESP_DLY3~q ),
	.prn(vcc));
defparam \ctrl_state.PUTRESP_DLY3 .is_wysiwyg = "true";
defparam \ctrl_state.PUTRESP_DLY3 .power_up = "low";

fiftyfivenm_lcell_comb \Selector6~1 (
	.dataa(\ctrl_state.WAIT~q ),
	.datab(\ctrl_state.PUTRESP_DLY3~q ),
	.datac(gnd),
	.datad(\pend~q ),
	.cin(gnd),
	.combout(\Selector6~1_combout ),
	.cout());
defparam \Selector6~1 .lut_mask = 16'hEEFF;
defparam \Selector6~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector6~2 (
	.dataa(\Selector6~1_combout ),
	.datab(gnd),
	.datac(\Selector7~0_combout ),
	.datad(cmd_eop),
	.cin(gnd),
	.combout(\Selector6~2_combout ),
	.cout());
defparam \Selector6~2 .lut_mask = 16'hAFFF;
defparam \Selector6~2 .sum_lutc_input = "datac";

dffeas \ctrl_state.WAIT (
	.clk(clk_clk),
	.d(\Selector6~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_state.WAIT~q ),
	.prn(vcc));
defparam \ctrl_state.WAIT .is_wysiwyg = "true";
defparam \ctrl_state.WAIT .power_up = "low";

fiftyfivenm_lcell_comb \ctrl_state_nxt.GETCMD_W~0 (
	.dataa(cmd_eop),
	.datab(\ctrl_state.WAIT~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\ctrl_state_nxt.GETCMD_W~0_combout ),
	.cout());
defparam \ctrl_state_nxt.GETCMD_W~0 .lut_mask = 16'hEEEE;
defparam \ctrl_state_nxt.GETCMD_W~0 .sum_lutc_input = "datac";

dffeas \ctrl_state.GETCMD_W (
	.clk(clk_clk),
	.d(\ctrl_state_nxt.GETCMD_W~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_state.GETCMD_W~q ),
	.prn(vcc));
defparam \ctrl_state.GETCMD_W .is_wysiwyg = "true";
defparam \ctrl_state.GETCMD_W .power_up = "low";

fiftyfivenm_lcell_comb \Selector1~0 (
	.dataa(cmd_channel_4),
	.datab(\ctrl_state.GETCMD_W~q ),
	.datac(\ctrl_state.GETCMD~q ),
	.datad(\pend~q ),
	.cin(gnd),
	.combout(\Selector1~0_combout ),
	.cout());
defparam \Selector1~0 .lut_mask = 16'hFEFF;
defparam \Selector1~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector1~2 (
	.dataa(\Selector1~0_combout ),
	.datab(\Selector1~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector1~2_combout ),
	.cout());
defparam \Selector1~2 .lut_mask = 16'hEEEE;
defparam \Selector1~2 .sum_lutc_input = "datac";

dffeas \ctrl_state.PWRDWN (
	.clk(clk_clk),
	.d(\Selector1~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_state.PWRDWN~q ),
	.prn(vcc));
defparam \ctrl_state.PWRDWN .is_wysiwyg = "true";
defparam \ctrl_state.PWRDWN .power_up = "low";

fiftyfivenm_lcell_comb \Add0~0 (
	.dataa(\int_timer[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout(\Add0~1 ));
defparam \Add0~0 .lut_mask = 16'h55AA;
defparam \Add0~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \int_timer~7 (
	.dataa(\Add0~0_combout ),
	.datab(\ctrl_state.CONV~q ),
	.datac(\Selector9~1_combout ),
	.datad(\cmd_fetched~0_combout ),
	.cin(gnd),
	.combout(\int_timer~7_combout ),
	.cout());
defparam \int_timer~7 .lut_mask = 16'hEFFF;
defparam \int_timer~7 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \load_int_timer~0 (
	.dataa(\cmd_fetched~0_combout ),
	.datab(\Selector9~1_combout ),
	.datac(gnd),
	.datad(\ctrl_state.CONV~q ),
	.cin(gnd),
	.combout(\load_int_timer~0_combout ),
	.cout());
defparam \load_int_timer~0 .lut_mask = 16'hEEFF;
defparam \load_int_timer~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add0~12 (
	.dataa(\int_timer[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~11 ),
	.combout(\Add0~12_combout ),
	.cout(\Add0~13 ));
defparam \Add0~12 .lut_mask = 16'h5AAF;
defparam \Add0~12 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add0~14 (
	.dataa(\int_timer[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add0~13 ),
	.combout(\Add0~14_combout ),
	.cout());
defparam \Add0~14 .lut_mask = 16'h5A5A;
defparam \Add0~14 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \int_timer~8 (
	.dataa(\Add0~14_combout ),
	.datab(\ctrl_state.CONV~q ),
	.datac(\Selector9~1_combout ),
	.datad(\cmd_fetched~0_combout ),
	.cin(gnd),
	.combout(\int_timer~8_combout ),
	.cout());
defparam \int_timer~8 .lut_mask = 16'hEFFF;
defparam \int_timer~8 .sum_lutc_input = "datac";

dffeas \int_timer[7] (
	.clk(clk_clk),
	.d(\int_timer~8_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\int_timer[6]~0_combout ),
	.q(\int_timer[7]~q ),
	.prn(vcc));
defparam \int_timer[7] .is_wysiwyg = "true";
defparam \int_timer[7] .power_up = "low";

fiftyfivenm_lcell_comb \Selector2~0 (
	.dataa(\int_timer[6]~q ),
	.datab(\ctrl_state.PWRDWN~q ),
	.datac(\ctrl_state.PWRDWN_TSEN~q ),
	.datad(\int_timer[7]~q ),
	.cin(gnd),
	.combout(\Selector2~0_combout ),
	.cout());
defparam \Selector2~0 .lut_mask = 16'hFEFF;
defparam \Selector2~0 .sum_lutc_input = "datac";

dffeas \ctrl_state.PWRDWN_TSEN (
	.clk(clk_clk),
	.d(\Selector2~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_state.PWRDWN_TSEN~q ),
	.prn(vcc));
defparam \ctrl_state.PWRDWN_TSEN .is_wysiwyg = "true";
defparam \ctrl_state.PWRDWN_TSEN .power_up = "low";

fiftyfivenm_lcell_comb \int_timer[6]~0 (
	.dataa(\ctrl_state.PWRDWN~q ),
	.datab(\load_int_timer~0_combout ),
	.datac(\ctrl_state.PWRDWN_TSEN~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\int_timer[6]~0_combout ),
	.cout());
defparam \int_timer[6]~0 .lut_mask = 16'hFEFE;
defparam \int_timer[6]~0 .sum_lutc_input = "datac";

dffeas \int_timer[0] (
	.clk(clk_clk),
	.d(\int_timer~7_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\int_timer[6]~0_combout ),
	.q(\int_timer[0]~q ),
	.prn(vcc));
defparam \int_timer[0] .is_wysiwyg = "true";
defparam \int_timer[0] .power_up = "low";

fiftyfivenm_lcell_comb \Add0~2 (
	.dataa(\int_timer[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~1 ),
	.combout(\Add0~2_combout ),
	.cout(\Add0~3 ));
defparam \Add0~2 .lut_mask = 16'h5A5F;
defparam \Add0~2 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \int_timer~6 (
	.dataa(\Add0~2_combout ),
	.datab(\ctrl_state.CONV~q ),
	.datac(\Selector9~1_combout ),
	.datad(\cmd_fetched~0_combout ),
	.cin(gnd),
	.combout(\int_timer~6_combout ),
	.cout());
defparam \int_timer~6 .lut_mask = 16'hEFFF;
defparam \int_timer~6 .sum_lutc_input = "datac";

dffeas \int_timer[1] (
	.clk(clk_clk),
	.d(\int_timer~6_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\int_timer[6]~0_combout ),
	.q(\int_timer[1]~q ),
	.prn(vcc));
defparam \int_timer[1] .is_wysiwyg = "true";
defparam \int_timer[1] .power_up = "low";

fiftyfivenm_lcell_comb \Add0~4 (
	.dataa(\int_timer[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~3 ),
	.combout(\Add0~4_combout ),
	.cout(\Add0~5 ));
defparam \Add0~4 .lut_mask = 16'h5AAF;
defparam \Add0~4 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \int_timer~5 (
	.dataa(\Add0~4_combout ),
	.datab(\ctrl_state.CONV~q ),
	.datac(\Selector9~1_combout ),
	.datad(\cmd_fetched~0_combout ),
	.cin(gnd),
	.combout(\int_timer~5_combout ),
	.cout());
defparam \int_timer~5 .lut_mask = 16'hEFFF;
defparam \int_timer~5 .sum_lutc_input = "datac";

dffeas \int_timer[2] (
	.clk(clk_clk),
	.d(\int_timer~5_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\int_timer[6]~0_combout ),
	.q(\int_timer[2]~q ),
	.prn(vcc));
defparam \int_timer[2] .is_wysiwyg = "true";
defparam \int_timer[2] .power_up = "low";

fiftyfivenm_lcell_comb \Add0~6 (
	.dataa(\int_timer[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~5 ),
	.combout(\Add0~6_combout ),
	.cout(\Add0~7 ));
defparam \Add0~6 .lut_mask = 16'h5A5F;
defparam \Add0~6 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \int_timer~4 (
	.dataa(\Add0~6_combout ),
	.datab(\ctrl_state.CONV~q ),
	.datac(\Selector9~1_combout ),
	.datad(\cmd_fetched~0_combout ),
	.cin(gnd),
	.combout(\int_timer~4_combout ),
	.cout());
defparam \int_timer~4 .lut_mask = 16'hEFFF;
defparam \int_timer~4 .sum_lutc_input = "datac";

dffeas \int_timer[3] (
	.clk(clk_clk),
	.d(\int_timer~4_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\int_timer[6]~0_combout ),
	.q(\int_timer[3]~q ),
	.prn(vcc));
defparam \int_timer[3] .is_wysiwyg = "true";
defparam \int_timer[3] .power_up = "low";

fiftyfivenm_lcell_comb \Add0~8 (
	.dataa(\int_timer[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~7 ),
	.combout(\Add0~8_combout ),
	.cout(\Add0~9 ));
defparam \Add0~8 .lut_mask = 16'h5AAF;
defparam \Add0~8 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \int_timer~3 (
	.dataa(\Add0~8_combout ),
	.datab(\ctrl_state.CONV~q ),
	.datac(\Selector9~1_combout ),
	.datad(\cmd_fetched~0_combout ),
	.cin(gnd),
	.combout(\int_timer~3_combout ),
	.cout());
defparam \int_timer~3 .lut_mask = 16'hEFFF;
defparam \int_timer~3 .sum_lutc_input = "datac";

dffeas \int_timer[4] (
	.clk(clk_clk),
	.d(\int_timer~3_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\int_timer[6]~0_combout ),
	.q(\int_timer[4]~q ),
	.prn(vcc));
defparam \int_timer[4] .is_wysiwyg = "true";
defparam \int_timer[4] .power_up = "low";

fiftyfivenm_lcell_comb \Add0~10 (
	.dataa(\int_timer[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~9 ),
	.combout(\Add0~10_combout ),
	.cout(\Add0~11 ));
defparam \Add0~10 .lut_mask = 16'h5A5F;
defparam \Add0~10 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \int_timer~2 (
	.dataa(\Add0~10_combout ),
	.datab(\ctrl_state.CONV~q ),
	.datac(\Selector9~1_combout ),
	.datad(\cmd_fetched~0_combout ),
	.cin(gnd),
	.combout(\int_timer~2_combout ),
	.cout());
defparam \int_timer~2 .lut_mask = 16'hEFFF;
defparam \int_timer~2 .sum_lutc_input = "datac";

dffeas \int_timer[5] (
	.clk(clk_clk),
	.d(\int_timer~2_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\int_timer[6]~0_combout ),
	.q(\int_timer[5]~q ),
	.prn(vcc));
defparam \int_timer[5] .is_wysiwyg = "true";
defparam \int_timer[5] .power_up = "low";

fiftyfivenm_lcell_comb \int_timer[6]~1 (
	.dataa(\int_timer[6]~q ),
	.datab(\Add0~12_combout ),
	.datac(\int_timer[6]~0_combout ),
	.datad(\load_int_timer~0_combout ),
	.cin(gnd),
	.combout(\int_timer[6]~1_combout ),
	.cout());
defparam \int_timer[6]~1 .lut_mask = 16'hACFF;
defparam \int_timer[6]~1 .sum_lutc_input = "datac";

dffeas \int_timer[6] (
	.clk(clk_clk),
	.d(\int_timer[6]~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\int_timer[6]~q ),
	.prn(vcc));
defparam \int_timer[6] .is_wysiwyg = "true";
defparam \int_timer[6] .power_up = "low";

fiftyfivenm_lcell_comb \Selector0~0 (
	.dataa(wire_pll7_locked),
	.datab(\ctrl_state.IDLE~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector0~0_combout ),
	.cout());
defparam \Selector0~0 .lut_mask = 16'hEEEE;
defparam \Selector0~0 .sum_lutc_input = "datac";

dffeas \ctrl_state.IDLE (
	.clk(clk_clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_state.IDLE~q ),
	.prn(vcc));
defparam \ctrl_state.IDLE .is_wysiwyg = "true";
defparam \ctrl_state.IDLE .power_up = "low";

fiftyfivenm_lcell_comb \Selector1~1 (
	.dataa(\ctrl_state.PWRDWN~q ),
	.datab(wire_pll7_locked),
	.datac(\int_timer[6]~q ),
	.datad(\ctrl_state.IDLE~q ),
	.cin(gnd),
	.combout(\Selector1~1_combout ),
	.cout());
defparam \Selector1~1 .lut_mask = 16'hEFFF;
defparam \Selector1~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \cmd_fetched~0 (
	.dataa(\ctrl_state.GETCMD~q ),
	.datab(\ctrl_state.GETCMD_W~q ),
	.datac(\Selector1~0_combout ),
	.datad(\Selector1~1_combout ),
	.cin(gnd),
	.combout(\cmd_fetched~0_combout ),
	.cout());
defparam \cmd_fetched~0 .lut_mask = 16'hFFFE;
defparam \cmd_fetched~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector5~0 (
	.dataa(\ctrl_state.PWRUP_SOC~q ),
	.datab(\u_eoc_synchronizer|dreg[0]~q ),
	.datac(gnd),
	.datad(\eoc_synch_dly~q ),
	.cin(gnd),
	.combout(\Selector5~0_combout ),
	.cout());
defparam \Selector5~0 .lut_mask = 16'hEEFF;
defparam \Selector5~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector3~0 (
	.dataa(\ctrl_state.PWRDWN_TSEN~q ),
	.datab(\int_timer[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector3~0_combout ),
	.cout());
defparam \Selector3~0 .lut_mask = 16'hEEEE;
defparam \Selector3~0 .sum_lutc_input = "datac";

dffeas clk_dft_synch_dly(
	.clk(clk_clk),
	.d(\u_clk_dft_synchronizer|dreg[0]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\clk_dft_synch_dly~q ),
	.prn(vcc));
defparam clk_dft_synch_dly.is_wysiwyg = "true";
defparam clk_dft_synch_dly.power_up = "low";

fiftyfivenm_lcell_comb \Selector3~1 (
	.dataa(\Selector3~0_combout ),
	.datab(\ctrl_state.PWRDWN_DONE~q ),
	.datac(\clk_dft_synch_dly~q ),
	.datad(\u_clk_dft_synchronizer|dreg[0]~q ),
	.cin(gnd),
	.combout(\Selector3~1_combout ),
	.cout());
defparam \Selector3~1 .lut_mask = 16'hFEFF;
defparam \Selector3~1 .sum_lutc_input = "datac";

dffeas \ctrl_state.PWRDWN_DONE (
	.clk(clk_clk),
	.d(\Selector3~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_state.PWRDWN_DONE~q ),
	.prn(vcc));
defparam \ctrl_state.PWRDWN_DONE .is_wysiwyg = "true";
defparam \ctrl_state.PWRDWN_DONE .power_up = "low";

fiftyfivenm_lcell_comb \Selector4~0 (
	.dataa(\ctrl_state.PWRUP_CH~q ),
	.datab(\u_clk_dft_synchronizer|dreg[0]~q ),
	.datac(\ctrl_state.PWRDWN_DONE~q ),
	.datad(\clk_dft_synch_dly~q ),
	.cin(gnd),
	.combout(\Selector4~0_combout ),
	.cout());
defparam \Selector4~0 .lut_mask = 16'hFEFF;
defparam \Selector4~0 .sum_lutc_input = "datac";

dffeas \ctrl_state.PWRUP_CH (
	.clk(clk_clk),
	.d(\Selector4~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_state.PWRUP_CH~q ),
	.prn(vcc));
defparam \ctrl_state.PWRUP_CH .is_wysiwyg = "true";
defparam \ctrl_state.PWRUP_CH .power_up = "low";

fiftyfivenm_lcell_comb \Selector5~1 (
	.dataa(\Selector5~0_combout ),
	.datab(\ctrl_state.PWRUP_CH~q ),
	.datac(\clk_dft_synch_dly~q ),
	.datad(\u_clk_dft_synchronizer|dreg[0]~q ),
	.cin(gnd),
	.combout(\Selector5~1_combout ),
	.cout());
defparam \Selector5~1 .lut_mask = 16'hFEFF;
defparam \Selector5~1 .sum_lutc_input = "datac";

dffeas \ctrl_state.PWRUP_SOC (
	.clk(clk_clk),
	.d(\Selector5~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_state.PWRUP_SOC~q ),
	.prn(vcc));
defparam \ctrl_state.PWRUP_SOC .is_wysiwyg = "true";
defparam \ctrl_state.PWRUP_SOC .power_up = "low";

fiftyfivenm_lcell_comb \Selector6~0 (
	.dataa(\ctrl_state.PWRUP_SOC~q ),
	.datab(\eoc_synch_dly~q ),
	.datac(gnd),
	.datad(\u_eoc_synchronizer|dreg[0]~q ),
	.cin(gnd),
	.combout(\Selector6~0_combout ),
	.cout());
defparam \Selector6~0 .lut_mask = 16'hEEFF;
defparam \Selector6~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \cmd_fetched~1 (
	.dataa(\cmd_fetched~0_combout ),
	.datab(\cmd_fetched~q ),
	.datac(gnd),
	.datad(\Selector6~0_combout ),
	.cin(gnd),
	.combout(\cmd_fetched~1_combout ),
	.cout());
defparam \cmd_fetched~1 .lut_mask = 16'hEEFF;
defparam \cmd_fetched~1 .sum_lutc_input = "datac";

dffeas cmd_fetched(
	.clk(clk_clk),
	.d(\cmd_fetched~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\cmd_fetched~q ),
	.prn(vcc));
defparam cmd_fetched.is_wysiwyg = "true";
defparam cmd_fetched.power_up = "low";

fiftyfivenm_lcell_comb \Selector7~0 (
	.dataa(\cmd_fetched~q ),
	.datab(gnd),
	.datac(\Selector6~0_combout ),
	.datad(\ctrl_state.PUTRESP_PEND~q ),
	.cin(gnd),
	.combout(\Selector7~0_combout ),
	.cout());
defparam \Selector7~0 .lut_mask = 16'hAFFF;
defparam \Selector7~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector7~1 (
	.dataa(cmd_eop),
	.datab(\ctrl_state.PUTRESP_DLY3~q ),
	.datac(gnd),
	.datad(\Selector7~0_combout ),
	.cin(gnd),
	.combout(\Selector7~1_combout ),
	.cout());
defparam \Selector7~1 .lut_mask = 16'hEEFF;
defparam \Selector7~1 .sum_lutc_input = "datac";

dffeas \ctrl_state.GETCMD (
	.clk(clk_clk),
	.d(\Selector7~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_state.GETCMD~q ),
	.prn(vcc));
defparam \ctrl_state.GETCMD .is_wysiwyg = "true";
defparam \ctrl_state.GETCMD .power_up = "low";

fiftyfivenm_lcell_comb \Selector9~0 (
	.dataa(\ctrl_state.GETCMD~q ),
	.datab(\cmd_fetched~q ),
	.datac(\Selector6~0_combout ),
	.datad(cmd_channel_4),
	.cin(gnd),
	.combout(\Selector9~0_combout ),
	.cout());
defparam \Selector9~0 .lut_mask = 16'hFEFF;
defparam \Selector9~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \ctrl_state_nxt~0 (
	.dataa(\eoc_synch_dly~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\u_eoc_synchronizer|dreg[0]~q ),
	.cin(gnd),
	.combout(\ctrl_state_nxt~0_combout ),
	.cout());
defparam \ctrl_state_nxt~0 .lut_mask = 16'hAAFF;
defparam \ctrl_state_nxt~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector8~0 (
	.dataa(\ctrl_state.GETCMD_W~q ),
	.datab(\ctrl_state.PRE_CONV~q ),
	.datac(cmd_channel_4),
	.datad(\ctrl_state_nxt~0_combout ),
	.cin(gnd),
	.combout(\Selector8~0_combout ),
	.cout());
defparam \Selector8~0 .lut_mask = 16'hEFFF;
defparam \Selector8~0 .sum_lutc_input = "datac";

dffeas \ctrl_state.PRE_CONV (
	.clk(clk_clk),
	.d(\Selector8~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_state.PRE_CONV~q ),
	.prn(vcc));
defparam \ctrl_state.PRE_CONV .is_wysiwyg = "true";
defparam \ctrl_state.PRE_CONV .power_up = "low";

fiftyfivenm_lcell_comb \Selector9~1 (
	.dataa(\Selector9~0_combout ),
	.datab(\ctrl_state.PRE_CONV~q ),
	.datac(\ctrl_state.CONV~q ),
	.datad(\ctrl_state_nxt~0_combout ),
	.cin(gnd),
	.combout(\Selector9~1_combout ),
	.cout());
defparam \Selector9~1 .lut_mask = 16'hFAFC;
defparam \Selector9~1 .sum_lutc_input = "datac";

dffeas \ctrl_state.CONV (
	.clk(clk_clk),
	.d(\Selector9~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_state.CONV~q ),
	.prn(vcc));
defparam \ctrl_state.CONV .is_wysiwyg = "true";
defparam \ctrl_state.CONV .power_up = "low";

fiftyfivenm_lcell_comb \ctrl_state_nxt.CONV_DLY1~0 (
	.dataa(\eoc_synch_dly~q ),
	.datab(\ctrl_state.CONV~q ),
	.datac(gnd),
	.datad(\u_eoc_synchronizer|dreg[0]~q ),
	.cin(gnd),
	.combout(\ctrl_state_nxt.CONV_DLY1~0_combout ),
	.cout());
defparam \ctrl_state_nxt.CONV_DLY1~0 .lut_mask = 16'hEEFF;
defparam \ctrl_state_nxt.CONV_DLY1~0 .sum_lutc_input = "datac";

dffeas \ctrl_state.CONV_DLY1 (
	.clk(clk_clk),
	.d(\ctrl_state_nxt.CONV_DLY1~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_state.CONV_DLY1~q ),
	.prn(vcc));
defparam \ctrl_state.CONV_DLY1 .is_wysiwyg = "true";
defparam \ctrl_state.CONV_DLY1 .power_up = "low";

dffeas conv_dly1_s_flp(
	.clk(clk_clk),
	.d(\ctrl_state.CONV_DLY1~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\conv_dly1_s_flp~q ),
	.prn(vcc));
defparam conv_dly1_s_flp.is_wysiwyg = "true";
defparam conv_dly1_s_flp.power_up = "low";

fiftyfivenm_lcell_comb \pend~0 (
	.dataa(\conv_dly1_s_flp~q ),
	.datab(\pend~q ),
	.datac(gnd),
	.datad(\ctrl_state.WAIT_PEND_DLY1~q ),
	.cin(gnd),
	.combout(\pend~0_combout ),
	.cout());
defparam \pend~0 .lut_mask = 16'hEEFF;
defparam \pend~0 .sum_lutc_input = "datac";

dffeas pend(
	.clk(clk_clk),
	.d(\pend~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pend~q ),
	.prn(vcc));
defparam pend.is_wysiwyg = "true";
defparam pend.power_up = "low";

fiftyfivenm_lcell_comb \Selector11~0 (
	.dataa(cmd_channel_4),
	.datab(\ctrl_state.GETCMD~q ),
	.datac(\ctrl_state.PUTRESP_DLY3~q ),
	.datad(cmd_eop),
	.cin(gnd),
	.combout(\Selector11~0_combout ),
	.cout());
defparam \Selector11~0 .lut_mask = 16'hFEFF;
defparam \Selector11~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector11~1 (
	.dataa(\pend~q ),
	.datab(\Selector11~0_combout ),
	.datac(\ctrl_state.WAIT_PEND~q ),
	.datad(\ctrl_state_nxt~0_combout ),
	.cin(gnd),
	.combout(\Selector11~1_combout ),
	.cout());
defparam \Selector11~1 .lut_mask = 16'hFEFF;
defparam \Selector11~1 .sum_lutc_input = "datac";

dffeas \ctrl_state.WAIT_PEND (
	.clk(clk_clk),
	.d(\Selector11~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_state.WAIT_PEND~q ),
	.prn(vcc));
defparam \ctrl_state.WAIT_PEND .is_wysiwyg = "true";
defparam \ctrl_state.WAIT_PEND .power_up = "low";

fiftyfivenm_lcell_comb \ctrl_state_nxt.WAIT_PEND_DLY1~0 (
	.dataa(\eoc_synch_dly~q ),
	.datab(\ctrl_state.WAIT_PEND~q ),
	.datac(gnd),
	.datad(\u_eoc_synchronizer|dreg[0]~q ),
	.cin(gnd),
	.combout(\ctrl_state_nxt.WAIT_PEND_DLY1~0_combout ),
	.cout());
defparam \ctrl_state_nxt.WAIT_PEND_DLY1~0 .lut_mask = 16'hEEFF;
defparam \ctrl_state_nxt.WAIT_PEND_DLY1~0 .sum_lutc_input = "datac";

dffeas \ctrl_state.WAIT_PEND_DLY1 (
	.clk(clk_clk),
	.d(\ctrl_state_nxt.WAIT_PEND_DLY1~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_state.WAIT_PEND_DLY1~q ),
	.prn(vcc));
defparam \ctrl_state.WAIT_PEND_DLY1 .is_wysiwyg = "true";
defparam \ctrl_state.WAIT_PEND_DLY1 .power_up = "low";

dffeas \ctrl_state.PUTRESP_PEND (
	.clk(clk_clk),
	.d(\ctrl_state.WAIT_PEND_DLY1~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_state.PUTRESP_PEND~q ),
	.prn(vcc));
defparam \ctrl_state.PUTRESP_PEND .is_wysiwyg = "true";
defparam \ctrl_state.PUTRESP_PEND .power_up = "low";

fiftyfivenm_lcell_comb \Selector10~0 (
	.dataa(\ctrl_state.CONV_DLY1~q ),
	.datab(cmd_channel_4),
	.datac(\cmd_fetched~q ),
	.datad(\Selector6~0_combout ),
	.cin(gnd),
	.combout(\Selector10~0_combout ),
	.cout());
defparam \Selector10~0 .lut_mask = 16'hFFFE;
defparam \Selector10~0 .sum_lutc_input = "datac";

dffeas \ctrl_state.PUTRESP (
	.clk(clk_clk),
	.d(\Selector10~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ctrl_state.PUTRESP~q ),
	.prn(vcc));
defparam \ctrl_state.PUTRESP .is_wysiwyg = "true";
defparam \ctrl_state.PUTRESP .power_up = "low";

fiftyfivenm_lcell_comb load_rsp(
	.dataa(\ctrl_state.PUTRESP_PEND~q ),
	.datab(\ctrl_state.PUTRESP~q ),
	.datac(\pend~q ),
	.datad(cmd_channel_4),
	.cin(gnd),
	.combout(\load_rsp~combout ),
	.cout());
defparam load_rsp.lut_mask = 16'hFEFF;
defparam load_rsp.sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \load_dout~2 (
	.dataa(\ctrl_state.WAIT_PEND~q ),
	.datab(\pend~q ),
	.datac(\ctrl_state.CONV~q ),
	.datad(cmd_channel_4),
	.cin(gnd),
	.combout(\load_dout~2_combout ),
	.cout());
defparam \load_dout~2 .lut_mask = 16'hFEFF;
defparam \load_dout~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \load_dout~3 (
	.dataa(\eoc_synch_dly~q ),
	.datab(\u_eoc_synchronizer|dreg[0]~q ),
	.datac(\load_dout~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\load_dout~3_combout ),
	.cout());
defparam \load_dout~3 .lut_mask = 16'hFBFB;
defparam \load_dout~3 .sum_lutc_input = "datac";

dffeas \dout_flp[0] (
	.clk(clk_clk),
	.d(wire_from_adc_dout_0),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_dout~3_combout ),
	.q(\dout_flp[0]~q ),
	.prn(vcc));
defparam \dout_flp[0] .is_wysiwyg = "true";
defparam \dout_flp[0] .power_up = "low";

fiftyfivenm_lcell_comb \rsp_data~0 (
	.dataa(\load_rsp~combout ),
	.datab(\dout_flp[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rsp_data~0_combout ),
	.cout());
defparam \rsp_data~0 .lut_mask = 16'hEEEE;
defparam \rsp_data~0 .sum_lutc_input = "datac";

dffeas \dout_flp[2] (
	.clk(clk_clk),
	.d(wire_from_adc_dout_2),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_dout~3_combout ),
	.q(\dout_flp[2]~q ),
	.prn(vcc));
defparam \dout_flp[2] .is_wysiwyg = "true";
defparam \dout_flp[2] .power_up = "low";

fiftyfivenm_lcell_comb \rsp_data~1 (
	.dataa(\load_rsp~combout ),
	.datab(\dout_flp[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rsp_data~1_combout ),
	.cout());
defparam \rsp_data~1 .lut_mask = 16'hEEEE;
defparam \rsp_data~1 .sum_lutc_input = "datac";

dffeas \dout_flp[1] (
	.clk(clk_clk),
	.d(wire_from_adc_dout_1),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_dout~3_combout ),
	.q(\dout_flp[1]~q ),
	.prn(vcc));
defparam \dout_flp[1] .is_wysiwyg = "true";
defparam \dout_flp[1] .power_up = "low";

fiftyfivenm_lcell_comb \rsp_data~2 (
	.dataa(\load_rsp~combout ),
	.datab(\dout_flp[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rsp_data~2_combout ),
	.cout());
defparam \rsp_data~2 .lut_mask = 16'hEEEE;
defparam \rsp_data~2 .sum_lutc_input = "datac";

dffeas \dout_flp[5] (
	.clk(clk_clk),
	.d(wire_from_adc_dout_5),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_dout~3_combout ),
	.q(\dout_flp[5]~q ),
	.prn(vcc));
defparam \dout_flp[5] .is_wysiwyg = "true";
defparam \dout_flp[5] .power_up = "low";

fiftyfivenm_lcell_comb \rsp_data~3 (
	.dataa(\load_rsp~combout ),
	.datab(\dout_flp[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rsp_data~3_combout ),
	.cout());
defparam \rsp_data~3 .lut_mask = 16'hEEEE;
defparam \rsp_data~3 .sum_lutc_input = "datac";

dffeas \dout_flp[7] (
	.clk(clk_clk),
	.d(wire_from_adc_dout_7),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_dout~3_combout ),
	.q(\dout_flp[7]~q ),
	.prn(vcc));
defparam \dout_flp[7] .is_wysiwyg = "true";
defparam \dout_flp[7] .power_up = "low";

fiftyfivenm_lcell_comb \rsp_data~4 (
	.dataa(\load_rsp~combout ),
	.datab(\dout_flp[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rsp_data~4_combout ),
	.cout());
defparam \rsp_data~4 .lut_mask = 16'hEEEE;
defparam \rsp_data~4 .sum_lutc_input = "datac";

dffeas \dout_flp[6] (
	.clk(clk_clk),
	.d(wire_from_adc_dout_6),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_dout~3_combout ),
	.q(\dout_flp[6]~q ),
	.prn(vcc));
defparam \dout_flp[6] .is_wysiwyg = "true";
defparam \dout_flp[6] .power_up = "low";

fiftyfivenm_lcell_comb \rsp_data~5 (
	.dataa(\load_rsp~combout ),
	.datab(\dout_flp[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rsp_data~5_combout ),
	.cout());
defparam \rsp_data~5 .lut_mask = 16'hEEEE;
defparam \rsp_data~5 .sum_lutc_input = "datac";

dffeas \dout_flp[4] (
	.clk(clk_clk),
	.d(wire_from_adc_dout_4),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_dout~3_combout ),
	.q(\dout_flp[4]~q ),
	.prn(vcc));
defparam \dout_flp[4] .is_wysiwyg = "true";
defparam \dout_flp[4] .power_up = "low";

fiftyfivenm_lcell_comb \rsp_data~6 (
	.dataa(\load_rsp~combout ),
	.datab(\dout_flp[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rsp_data~6_combout ),
	.cout());
defparam \rsp_data~6 .lut_mask = 16'hEEEE;
defparam \rsp_data~6 .sum_lutc_input = "datac";

dffeas \dout_flp[3] (
	.clk(clk_clk),
	.d(wire_from_adc_dout_3),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_dout~3_combout ),
	.q(\dout_flp[3]~q ),
	.prn(vcc));
defparam \dout_flp[3] .is_wysiwyg = "true";
defparam \dout_flp[3] .power_up = "low";

fiftyfivenm_lcell_comb \rsp_data~7 (
	.dataa(\load_rsp~combout ),
	.datab(\dout_flp[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rsp_data~7_combout ),
	.cout());
defparam \rsp_data~7 .lut_mask = 16'hEEEE;
defparam \rsp_data~7 .sum_lutc_input = "datac";

dffeas \dout_flp[8] (
	.clk(clk_clk),
	.d(wire_from_adc_dout_8),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_dout~3_combout ),
	.q(\dout_flp[8]~q ),
	.prn(vcc));
defparam \dout_flp[8] .is_wysiwyg = "true";
defparam \dout_flp[8] .power_up = "low";

fiftyfivenm_lcell_comb \rsp_data~8 (
	.dataa(\load_rsp~combout ),
	.datab(\dout_flp[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rsp_data~8_combout ),
	.cout());
defparam \rsp_data~8 .lut_mask = 16'hEEEE;
defparam \rsp_data~8 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \cmd_eop_dly~0 (
	.dataa(cmd_eop),
	.datab(\cmd_eop_dly~q ),
	.datac(gnd),
	.datad(\ctrl_state.PUTRESP~q ),
	.cin(gnd),
	.combout(\cmd_eop_dly~0_combout ),
	.cout());
defparam \cmd_eop_dly~0 .lut_mask = 16'hAACC;
defparam \cmd_eop_dly~0 .sum_lutc_input = "datac";

dffeas cmd_eop_dly(
	.clk(clk_clk),
	.d(\cmd_eop_dly~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\cmd_eop_dly~q ),
	.prn(vcc));
defparam cmd_eop_dly.is_wysiwyg = "true";
defparam cmd_eop_dly.power_up = "low";

fiftyfivenm_lcell_comb \rsp_eop~0 (
	.dataa(\load_rsp~combout ),
	.datab(\cmd_eop_dly~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rsp_eop~0_combout ),
	.cout());
defparam \rsp_eop~0 .lut_mask = 16'hEEEE;
defparam \rsp_eop~0 .sum_lutc_input = "datac";

dffeas \dout_flp[10] (
	.clk(clk_clk),
	.d(wire_from_adc_dout_10),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_dout~3_combout ),
	.q(\dout_flp[10]~q ),
	.prn(vcc));
defparam \dout_flp[10] .is_wysiwyg = "true";
defparam \dout_flp[10] .power_up = "low";

fiftyfivenm_lcell_comb \rsp_data~9 (
	.dataa(\load_rsp~combout ),
	.datab(\dout_flp[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rsp_data~9_combout ),
	.cout());
defparam \rsp_data~9 .lut_mask = 16'hEEEE;
defparam \rsp_data~9 .sum_lutc_input = "datac";

dffeas \dout_flp[9] (
	.clk(clk_clk),
	.d(wire_from_adc_dout_9),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_dout~3_combout ),
	.q(\dout_flp[9]~q ),
	.prn(vcc));
defparam \dout_flp[9] .is_wysiwyg = "true";
defparam \dout_flp[9] .power_up = "low";

fiftyfivenm_lcell_comb \rsp_data~10 (
	.dataa(\load_rsp~combout ),
	.datab(\dout_flp[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rsp_data~10_combout ),
	.cout());
defparam \rsp_data~10 .lut_mask = 16'hEEEE;
defparam \rsp_data~10 .sum_lutc_input = "datac";

dffeas \dout_flp[11] (
	.clk(clk_clk),
	.d(wire_from_adc_dout_11),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\load_dout~3_combout ),
	.q(\dout_flp[11]~q ),
	.prn(vcc));
defparam \dout_flp[11] .is_wysiwyg = "true";
defparam \dout_flp[11] .power_up = "low";

fiftyfivenm_lcell_comb \rsp_data~11 (
	.dataa(\load_rsp~combout ),
	.datab(\dout_flp[11]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\rsp_data~11_combout ),
	.cout());
defparam \rsp_data~11 .lut_mask = 16'hEEEE;
defparam \rsp_data~11 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \WideOr12~0 (
	.dataa(\Selector7~0_combout ),
	.datab(cmd_eop),
	.datac(\Selector6~1_combout ),
	.datad(\ctrl_state.PUTRESP_DLY3~q ),
	.cin(gnd),
	.combout(\WideOr12~0_combout ),
	.cout());
defparam \WideOr12~0 .lut_mask = 16'h8BFF;
defparam \WideOr12~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \WideOr12~1 (
	.dataa(\ctrl_state_nxt~0_combout ),
	.datab(\ctrl_state.WAIT_PEND~q ),
	.datac(cmd_ready1),
	.datad(\Selector10~0_combout ),
	.cin(gnd),
	.combout(\WideOr12~1_combout ),
	.cout());
defparam \WideOr12~1 .lut_mask = 16'h7FFF;
defparam \WideOr12~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \WideOr12~2 (
	.dataa(\ctrl_state.PUTRESP~q ),
	.datab(\ctrl_state.WAIT_PEND_DLY1~q ),
	.datac(\ctrl_state_nxt.GETCMD_W~0_combout ),
	.datad(\ctrl_state.PUTRESP_DLY2~q ),
	.cin(gnd),
	.combout(\WideOr12~2_combout ),
	.cout());
defparam \WideOr12~2 .lut_mask = 16'h7FFF;
defparam \WideOr12~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \WideOr12~3 (
	.dataa(\WideOr12~0_combout ),
	.datab(\WideOr12~1_combout ),
	.datac(\WideOr12~2_combout ),
	.datad(\Selector8~0_combout ),
	.cin(gnd),
	.combout(\WideOr12~3_combout ),
	.cout());
defparam \WideOr12~3 .lut_mask = 16'hFEFF;
defparam \WideOr12~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \WideOr13~0 (
	.dataa(\ctrl_state_nxt~0_combout ),
	.datab(\ctrl_state.PRE_CONV~q ),
	.datac(\ctrl_state.CONV~q ),
	.datad(\Selector9~0_combout ),
	.cin(gnd),
	.combout(\WideOr13~0_combout ),
	.cout());
defparam \WideOr13~0 .lut_mask = 16'h7FFF;
defparam \WideOr13~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \WideOr15~0 (
	.dataa(\WideOr12~3_combout ),
	.datab(\WideOr13~0_combout ),
	.datac(gnd),
	.datad(\Selector11~1_combout ),
	.cin(gnd),
	.combout(\WideOr15~0_combout ),
	.cout());
defparam \WideOr15~0 .lut_mask = 16'hEEFF;
defparam \WideOr15~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector17~0 (
	.dataa(\Selector5~1_combout ),
	.datab(soc1),
	.datac(\Selector4~0_combout ),
	.datad(\WideOr15~0_combout ),
	.cin(gnd),
	.combout(\Selector17~0_combout ),
	.cout());
defparam \Selector17~0 .lut_mask = 16'hFEFF;
defparam \Selector17~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \WideOr12~4 (
	.dataa(\Selector1~0_combout ),
	.datab(\Selector1~1_combout ),
	.datac(\Selector4~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\WideOr12~4_combout ),
	.cout());
defparam \WideOr12~4 .lut_mask = 16'hFEFE;
defparam \WideOr12~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb WideOr12(
	.dataa(\Selector5~1_combout ),
	.datab(\Selector3~1_combout ),
	.datac(\WideOr12~4_combout ),
	.datad(\WideOr12~3_combout ),
	.cin(gnd),
	.combout(\WideOr12~combout ),
	.cout());
defparam WideOr12.lut_mask = 16'hFEFF;
defparam WideOr12.sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector15~0 (
	.dataa(cmd_channel_4),
	.datab(\WideOr13~0_combout ),
	.datac(chsel_1),
	.datad(\WideOr12~combout ),
	.cin(gnd),
	.combout(\Selector15~0_combout ),
	.cout());
defparam \Selector15~0 .lut_mask = 16'hFFF7;
defparam \Selector15~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector16~0 (
	.dataa(chsel_0),
	.datab(\WideOr12~combout ),
	.datac(cmd_channel_4),
	.datad(\WideOr13~0_combout ),
	.cin(gnd),
	.combout(\Selector16~0_combout ),
	.cout());
defparam \Selector16~0 .lut_mask = 16'hFEFF;
defparam \Selector16~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector18~0 (
	.dataa(\Selector5~1_combout ),
	.datab(gnd),
	.datac(\WideOr15~0_combout ),
	.datad(\usr_pwd~q ),
	.cin(gnd),
	.combout(\Selector18~0_combout ),
	.cout());
defparam \Selector18~0 .lut_mask = 16'hAFFF;
defparam \Selector18~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector18~1 (
	.dataa(\Selector1~2_combout ),
	.datab(\Selector18~0_combout ),
	.datac(\Selector2~0_combout ),
	.datad(\Selector0~0_combout ),
	.cin(gnd),
	.combout(\Selector18~1_combout ),
	.cout());
defparam \Selector18~1 .lut_mask = 16'hFF7F;
defparam \Selector18~1 .sum_lutc_input = "datac";

dffeas usr_pwd(
	.clk(clk_clk),
	.d(\Selector18~1_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\usr_pwd~q ),
	.prn(vcc));
defparam usr_pwd.is_wysiwyg = "true";
defparam usr_pwd.power_up = "low";

endmodule

module ADC_altera_std_synchronizer (
	din,
	reset_n,
	dreg_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	din;
input 	reset_n;
output 	dreg_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module ADC_altera_std_synchronizer_1 (
	din,
	reset_n,
	dreg_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	din;
input 	reset_n;
output 	dreg_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module ADC_fiftyfivenm_adcblock_top_wrapper (
	eoc,
	clkout_adccore,
	wire_from_adc_dout_0,
	wire_from_adc_dout_1,
	wire_from_adc_dout_2,
	wire_from_adc_dout_3,
	wire_from_adc_dout_4,
	wire_from_adc_dout_5,
	wire_from_adc_dout_6,
	wire_from_adc_dout_7,
	wire_from_adc_dout_8,
	wire_from_adc_dout_9,
	wire_from_adc_dout_10,
	wire_from_adc_dout_11,
	wire_pll7_clk_0,
	soc,
	chsel_1,
	chsel_0,
	GND_port,
	chsel_11,
	usr_pwd)/* synthesis synthesis_greybox=1 */;
output 	eoc;
output 	clkout_adccore;
output 	wire_from_adc_dout_0;
output 	wire_from_adc_dout_1;
output 	wire_from_adc_dout_2;
output 	wire_from_adc_dout_3;
output 	wire_from_adc_dout_4;
output 	wire_from_adc_dout_5;
output 	wire_from_adc_dout_6;
output 	wire_from_adc_dout_7;
output 	wire_from_adc_dout_8;
output 	wire_from_adc_dout_9;
output 	wire_from_adc_dout_10;
output 	wire_from_adc_dout_11;
input 	wire_pll7_clk_0;
input 	soc;
input 	chsel_1;
input 	chsel_0;
input 	GND_port;
input 	chsel_11;
input 	usr_pwd;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \decoder|WideOr4~0_combout ;
wire \decoder|WideOr2~0_combout ;


ADC_fiftyfivenm_adcblock_primitive_wrapper adcblock_instance(
	.eoc(eoc),
	.clkout_adccore(clkout_adccore),
	.dout({wire_from_adc_dout_11,wire_from_adc_dout_10,wire_from_adc_dout_9,wire_from_adc_dout_8,wire_from_adc_dout_7,wire_from_adc_dout_6,wire_from_adc_dout_5,wire_from_adc_dout_4,wire_from_adc_dout_3,wire_from_adc_dout_2,wire_from_adc_dout_1,wire_from_adc_dout_0}),
	.clkin_from_pll_c0(wire_pll7_clk_0),
	.soc(soc),
	.chsel({chsel_11,chsel_11,\decoder|WideOr2~0_combout ,\decoder|WideOr4~0_combout ,\decoder|WideOr4~0_combout }),
	.tsen(GND_port),
	.usr_pwd(usr_pwd));

ADC_chsel_code_converter_sw_to_hw decoder(
	.chsel_1(chsel_1),
	.chsel_0(chsel_0),
	.WideOr4(\decoder|WideOr4~0_combout ),
	.WideOr2(\decoder|WideOr2~0_combout ));

endmodule

module ADC_chsel_code_converter_sw_to_hw (
	chsel_1,
	chsel_0,
	WideOr4,
	WideOr2)/* synthesis synthesis_greybox=1 */;
input 	chsel_1;
input 	chsel_0;
output 	WideOr4;
output 	WideOr2;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fiftyfivenm_lcell_comb \WideOr4~0 (
	.dataa(chsel_1),
	.datab(chsel_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(WideOr4),
	.cout());
defparam \WideOr4~0 .lut_mask = 16'h7777;
defparam \WideOr4~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \WideOr2~0 (
	.dataa(chsel_0),
	.datab(gnd),
	.datac(gnd),
	.datad(chsel_1),
	.cin(gnd),
	.combout(WideOr2),
	.cout());
defparam \WideOr2~0 .lut_mask = 16'hAAFF;
defparam \WideOr2~0 .sum_lutc_input = "datac";

endmodule

module ADC_fiftyfivenm_adcblock_primitive_wrapper (
	eoc,
	clkout_adccore,
	dout,
	clkin_from_pll_c0,
	soc,
	chsel,
	tsen,
	usr_pwd)/* synthesis synthesis_greybox=1 */;
output 	eoc;
output 	clkout_adccore;
output 	[11:0] dout;
input 	clkin_from_pll_c0;
input 	soc;
input 	[4:0] chsel;
input 	tsen;
input 	usr_pwd;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [11:0] primitive_instance_DOUT_bus;

assign dout[0] = primitive_instance_DOUT_bus[0];
assign dout[1] = primitive_instance_DOUT_bus[1];
assign dout[2] = primitive_instance_DOUT_bus[2];
assign dout[3] = primitive_instance_DOUT_bus[3];
assign dout[4] = primitive_instance_DOUT_bus[4];
assign dout[5] = primitive_instance_DOUT_bus[5];
assign dout[6] = primitive_instance_DOUT_bus[6];
assign dout[7] = primitive_instance_DOUT_bus[7];
assign dout[8] = primitive_instance_DOUT_bus[8];
assign dout[9] = primitive_instance_DOUT_bus[9];
assign dout[10] = primitive_instance_DOUT_bus[10];
assign dout[11] = primitive_instance_DOUT_bus[11];

fiftyfivenm_adcblock primitive_instance(
	.soc(soc),
	.usr_pwd(usr_pwd),
	.tsen(tsen),
	.clkin_from_pll_c0(clkin_from_pll_c0),
	.chsel({chsel[3],chsel[3],chsel[2],chsel[0],chsel[0]}),
	.eoc(eoc),
	.dout(primitive_instance_DOUT_bus));
defparam primitive_instance.analog_input_pin_mask = 0;
defparam primitive_instance.clkdiv = 2;
defparam primitive_instance.device_partname_fivechar_prefix = "10m50";
defparam primitive_instance.is_this_first_or_second_adc = 1;
defparam primitive_instance.prescalar = 0;
defparam primitive_instance.pwd = 0;
defparam primitive_instance.refsel = 1;
defparam primitive_instance.reserve_block = "false";
defparam primitive_instance.testbits = 66;
defparam primitive_instance.tsclkdiv = 1;
defparam primitive_instance.tsclksel = 1;

endmodule

module ADC_altera_modular_adc_sample_store (
	readdata_0,
	mem_used_2,
	address_7,
	address_6,
	address_5,
	address_4,
	Equal0,
	address_3,
	address_8,
	hold_waitrequest,
	write,
	readdata_2,
	readdata_1,
	readdata_5,
	readdata_7,
	readdata_6,
	readdata_4,
	readdata_3,
	readdata_8,
	rst_n,
	address_2,
	write1,
	readdata_10,
	readdata_9,
	readdata_13,
	readdata_15,
	readdata_14,
	readdata_12,
	readdata_11,
	rsp_valid,
	rsp_data_0,
	writedata_0,
	rsp_data_2,
	rsp_data_1,
	rsp_data_5,
	rsp_data_7,
	rsp_data_6,
	rsp_data_4,
	rsp_data_3,
	rsp_data_8,
	rsp_eop,
	rsp_data_10,
	rsp_data_9,
	rsp_data_11,
	GND_port,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	readdata_0;
input 	mem_used_2;
input 	address_7;
input 	address_6;
input 	address_5;
input 	address_4;
input 	Equal0;
input 	address_3;
input 	address_8;
input 	hold_waitrequest;
input 	write;
output 	readdata_2;
output 	readdata_1;
output 	readdata_5;
output 	readdata_7;
output 	readdata_6;
output 	readdata_4;
output 	readdata_3;
output 	readdata_8;
input 	rst_n;
input 	address_2;
input 	write1;
output 	readdata_10;
output 	readdata_9;
output 	readdata_13;
output 	readdata_15;
output 	readdata_14;
output 	readdata_12;
output 	readdata_11;
input 	rsp_valid;
input 	rsp_data_0;
input 	writedata_0;
input 	rsp_data_2;
input 	rsp_data_1;
input 	rsp_data_5;
input 	rsp_data_7;
input 	rsp_data_6;
input 	rsp_data_4;
input 	rsp_data_3;
input 	rsp_data_8;
input 	rsp_eop;
input 	rsp_data_10;
input 	rsp_data_9;
input 	rsp_data_11;
input 	GND_port;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \u_ss_ram|altsyncram_component|auto_generated|q_b[0] ;
wire \u_ss_ram|altsyncram_component|auto_generated|q_b[2] ;
wire \u_ss_ram|altsyncram_component|auto_generated|q_b[1] ;
wire \u_ss_ram|altsyncram_component|auto_generated|q_b[5] ;
wire \u_ss_ram|altsyncram_component|auto_generated|q_b[7] ;
wire \u_ss_ram|altsyncram_component|auto_generated|q_b[6] ;
wire \u_ss_ram|altsyncram_component|auto_generated|q_b[4] ;
wire \u_ss_ram|altsyncram_component|auto_generated|q_b[3] ;
wire \u_ss_ram|altsyncram_component|auto_generated|q_b[8] ;
wire \slot_num[0]~q ;
wire \slot_num[1]~q ;
wire \slot_num[2]~q ;
wire \slot_num[3]~q ;
wire \slot_num[4]~q ;
wire \slot_num[5]~q ;
wire \u_ss_ram|altsyncram_component|auto_generated|q_b[10] ;
wire \u_ss_ram|altsyncram_component|auto_generated|q_b[9] ;
wire \u_ss_ram|altsyncram_component|auto_generated|q_b[13] ;
wire \u_ss_ram|altsyncram_component|auto_generated|q_b[15] ;
wire \u_ss_ram|altsyncram_component|auto_generated|q_b[14] ;
wire \u_ss_ram|altsyncram_component|auto_generated|q_b[12] ;
wire \u_ss_ram|altsyncram_component|auto_generated|q_b[11] ;
wire \slot_num[0]~7 ;
wire \slot_num[0]~6_combout ;
wire \slot_num[1]~9 ;
wire \slot_num[1]~8_combout ;
wire \slot_num[2]~11 ;
wire \slot_num[2]~10_combout ;
wire \slot_num[3]~13 ;
wire \slot_num[3]~12_combout ;
wire \slot_num[4]~15 ;
wire \slot_num[4]~14_combout ;
wire \slot_num[5]~16_combout ;
wire \set_eop~combout ;
wire \csr_readdata_nxt[0]~1_combout ;
wire \ier_wr_en~0_combout ;
wire \always1~0_combout ;
wire \s_eop~0_combout ;
wire \s_eop~q ;
wire \e_eop~0_combout ;
wire \e_eop~q ;
wire \csr_readdata_nxt[0]~0_combout ;
wire \csr_readdata_nxt[0]~2_combout ;
wire \csr_readdata[0]~q ;
wire \ram_rd_en~combout ;
wire \ram_rd_en_flp~q ;
wire \readdata_nxt[0]~0_combout ;
wire \readdata_nxt[2]~1_combout ;
wire \readdata_nxt[1]~2_combout ;
wire \readdata_nxt[5]~3_combout ;
wire \readdata_nxt[7]~4_combout ;
wire \readdata_nxt[6]~5_combout ;
wire \readdata_nxt[4]~6_combout ;
wire \readdata_nxt[3]~7_combout ;
wire \readdata_nxt[8]~8_combout ;
wire \readdata_nxt[10]~9_combout ;
wire \readdata_nxt[9]~10_combout ;
wire \readdata_nxt[13]~11_combout ;
wire \readdata_nxt[15]~12_combout ;
wire \readdata_nxt[14]~13_combout ;
wire \readdata_nxt[12]~14_combout ;
wire \readdata_nxt[11]~15_combout ;


ADC_altera_modular_adc_sample_store_ram u_ss_ram(
	.q_b_0(\u_ss_ram|altsyncram_component|auto_generated|q_b[0] ),
	.q_b_2(\u_ss_ram|altsyncram_component|auto_generated|q_b[2] ),
	.q_b_1(\u_ss_ram|altsyncram_component|auto_generated|q_b[1] ),
	.q_b_5(\u_ss_ram|altsyncram_component|auto_generated|q_b[5] ),
	.q_b_7(\u_ss_ram|altsyncram_component|auto_generated|q_b[7] ),
	.q_b_6(\u_ss_ram|altsyncram_component|auto_generated|q_b[6] ),
	.q_b_4(\u_ss_ram|altsyncram_component|auto_generated|q_b[4] ),
	.q_b_3(\u_ss_ram|altsyncram_component|auto_generated|q_b[3] ),
	.q_b_8(\u_ss_ram|altsyncram_component|auto_generated|q_b[8] ),
	.slot_num_0(\slot_num[0]~q ),
	.slot_num_1(\slot_num[1]~q ),
	.slot_num_2(\slot_num[2]~q ),
	.slot_num_3(\slot_num[3]~q ),
	.slot_num_4(\slot_num[4]~q ),
	.slot_num_5(\slot_num[5]~q ),
	.q_b_10(\u_ss_ram|altsyncram_component|auto_generated|q_b[10] ),
	.q_b_9(\u_ss_ram|altsyncram_component|auto_generated|q_b[9] ),
	.q_b_13(\u_ss_ram|altsyncram_component|auto_generated|q_b[13] ),
	.q_b_15(\u_ss_ram|altsyncram_component|auto_generated|q_b[15] ),
	.q_b_14(\u_ss_ram|altsyncram_component|auto_generated|q_b[14] ),
	.q_b_12(\u_ss_ram|altsyncram_component|auto_generated|q_b[12] ),
	.q_b_11(\u_ss_ram|altsyncram_component|auto_generated|q_b[11] ),
	.address_7(address_7),
	.address_6(address_6),
	.address_5(address_5),
	.address_4(address_4),
	.address_3(address_3),
	.address_2(address_2),
	.rsp_valid(rsp_valid),
	.ram_rd_en(\ram_rd_en~combout ),
	.rsp_data_0(rsp_data_0),
	.rsp_data_2(rsp_data_2),
	.rsp_data_1(rsp_data_1),
	.rsp_data_5(rsp_data_5),
	.rsp_data_7(rsp_data_7),
	.rsp_data_6(rsp_data_6),
	.rsp_data_4(rsp_data_4),
	.rsp_data_3(rsp_data_3),
	.rsp_data_8(rsp_data_8),
	.rsp_data_10(rsp_data_10),
	.rsp_data_9(rsp_data_9),
	.rsp_data_11(rsp_data_11),
	.GND_port(GND_port),
	.clk_clk(clk_clk));

dffeas \slot_num[0] (
	.clk(clk_clk),
	.d(\slot_num[0]~6_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\set_eop~combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\slot_num[0]~q ),
	.prn(vcc));
defparam \slot_num[0] .is_wysiwyg = "true";
defparam \slot_num[0] .power_up = "low";

dffeas \slot_num[1] (
	.clk(clk_clk),
	.d(\slot_num[1]~8_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\set_eop~combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\slot_num[1]~q ),
	.prn(vcc));
defparam \slot_num[1] .is_wysiwyg = "true";
defparam \slot_num[1] .power_up = "low";

dffeas \slot_num[2] (
	.clk(clk_clk),
	.d(\slot_num[2]~10_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\set_eop~combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\slot_num[2]~q ),
	.prn(vcc));
defparam \slot_num[2] .is_wysiwyg = "true";
defparam \slot_num[2] .power_up = "low";

dffeas \slot_num[3] (
	.clk(clk_clk),
	.d(\slot_num[3]~12_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\set_eop~combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\slot_num[3]~q ),
	.prn(vcc));
defparam \slot_num[3] .is_wysiwyg = "true";
defparam \slot_num[3] .power_up = "low";

dffeas \slot_num[4] (
	.clk(clk_clk),
	.d(\slot_num[4]~14_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\set_eop~combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\slot_num[4]~q ),
	.prn(vcc));
defparam \slot_num[4] .is_wysiwyg = "true";
defparam \slot_num[4] .power_up = "low";

dffeas \slot_num[5] (
	.clk(clk_clk),
	.d(\slot_num[5]~16_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(\set_eop~combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\slot_num[5]~q ),
	.prn(vcc));
defparam \slot_num[5] .is_wysiwyg = "true";
defparam \slot_num[5] .power_up = "low";

fiftyfivenm_lcell_comb \slot_num[0]~6 (
	.dataa(\slot_num[0]~q ),
	.datab(rsp_valid),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\slot_num[0]~6_combout ),
	.cout(\slot_num[0]~7 ));
defparam \slot_num[0]~6 .lut_mask = 16'h66EE;
defparam \slot_num[0]~6 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \slot_num[1]~8 (
	.dataa(\slot_num[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\slot_num[0]~7 ),
	.combout(\slot_num[1]~8_combout ),
	.cout(\slot_num[1]~9 ));
defparam \slot_num[1]~8 .lut_mask = 16'h5A5F;
defparam \slot_num[1]~8 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \slot_num[2]~10 (
	.dataa(\slot_num[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\slot_num[1]~9 ),
	.combout(\slot_num[2]~10_combout ),
	.cout(\slot_num[2]~11 ));
defparam \slot_num[2]~10 .lut_mask = 16'h5AAF;
defparam \slot_num[2]~10 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \slot_num[3]~12 (
	.dataa(\slot_num[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\slot_num[2]~11 ),
	.combout(\slot_num[3]~12_combout ),
	.cout(\slot_num[3]~13 ));
defparam \slot_num[3]~12 .lut_mask = 16'h5A5F;
defparam \slot_num[3]~12 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \slot_num[4]~14 (
	.dataa(\slot_num[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\slot_num[3]~13 ),
	.combout(\slot_num[4]~14_combout ),
	.cout(\slot_num[4]~15 ));
defparam \slot_num[4]~14 .lut_mask = 16'h5AAF;
defparam \slot_num[4]~14 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \slot_num[5]~16 (
	.dataa(\slot_num[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\slot_num[4]~15 ),
	.combout(\slot_num[5]~16_combout ),
	.cout());
defparam \slot_num[5]~16 .lut_mask = 16'h5A5A;
defparam \slot_num[5]~16 .sum_lutc_input = "cin";

dffeas \readdata[0] (
	.clk(clk_clk),
	.d(\readdata_nxt[0]~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk_clk),
	.d(\readdata_nxt[2]~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk_clk),
	.d(\readdata_nxt[1]~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[5] (
	.clk(clk_clk),
	.d(\readdata_nxt[5]~3_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_5),
	.prn(vcc));
defparam \readdata[5] .is_wysiwyg = "true";
defparam \readdata[5] .power_up = "low";

dffeas \readdata[7] (
	.clk(clk_clk),
	.d(\readdata_nxt[7]~4_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_7),
	.prn(vcc));
defparam \readdata[7] .is_wysiwyg = "true";
defparam \readdata[7] .power_up = "low";

dffeas \readdata[6] (
	.clk(clk_clk),
	.d(\readdata_nxt[6]~5_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_6),
	.prn(vcc));
defparam \readdata[6] .is_wysiwyg = "true";
defparam \readdata[6] .power_up = "low";

dffeas \readdata[4] (
	.clk(clk_clk),
	.d(\readdata_nxt[4]~6_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_4),
	.prn(vcc));
defparam \readdata[4] .is_wysiwyg = "true";
defparam \readdata[4] .power_up = "low";

dffeas \readdata[3] (
	.clk(clk_clk),
	.d(\readdata_nxt[3]~7_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas \readdata[8] (
	.clk(clk_clk),
	.d(\readdata_nxt[8]~8_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_8),
	.prn(vcc));
defparam \readdata[8] .is_wysiwyg = "true";
defparam \readdata[8] .power_up = "low";

dffeas \readdata[10] (
	.clk(clk_clk),
	.d(\readdata_nxt[10]~9_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_10),
	.prn(vcc));
defparam \readdata[10] .is_wysiwyg = "true";
defparam \readdata[10] .power_up = "low";

dffeas \readdata[9] (
	.clk(clk_clk),
	.d(\readdata_nxt[9]~10_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_9),
	.prn(vcc));
defparam \readdata[9] .is_wysiwyg = "true";
defparam \readdata[9] .power_up = "low";

dffeas \readdata[13] (
	.clk(clk_clk),
	.d(\readdata_nxt[13]~11_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_13),
	.prn(vcc));
defparam \readdata[13] .is_wysiwyg = "true";
defparam \readdata[13] .power_up = "low";

dffeas \readdata[15] (
	.clk(clk_clk),
	.d(\readdata_nxt[15]~12_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_15),
	.prn(vcc));
defparam \readdata[15] .is_wysiwyg = "true";
defparam \readdata[15] .power_up = "low";

dffeas \readdata[14] (
	.clk(clk_clk),
	.d(\readdata_nxt[14]~13_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_14),
	.prn(vcc));
defparam \readdata[14] .is_wysiwyg = "true";
defparam \readdata[14] .power_up = "low";

dffeas \readdata[12] (
	.clk(clk_clk),
	.d(\readdata_nxt[12]~14_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_12),
	.prn(vcc));
defparam \readdata[12] .is_wysiwyg = "true";
defparam \readdata[12] .power_up = "low";

dffeas \readdata[11] (
	.clk(clk_clk),
	.d(\readdata_nxt[11]~15_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_11),
	.prn(vcc));
defparam \readdata[11] .is_wysiwyg = "true";
defparam \readdata[11] .power_up = "low";

fiftyfivenm_lcell_comb set_eop(
	.dataa(rsp_valid),
	.datab(rsp_eop),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\set_eop~combout ),
	.cout());
defparam set_eop.lut_mask = 16'hEEEE;
defparam set_eop.sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \csr_readdata_nxt[0]~1 (
	.dataa(Equal0),
	.datab(address_8),
	.datac(gnd),
	.datad(address_3),
	.cin(gnd),
	.combout(\csr_readdata_nxt[0]~1_combout ),
	.cout());
defparam \csr_readdata_nxt[0]~1 .lut_mask = 16'hEEFF;
defparam \csr_readdata_nxt[0]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \ier_wr_en~0 (
	.dataa(hold_waitrequest),
	.datab(write),
	.datac(\csr_readdata_nxt[0]~1_combout ),
	.datad(mem_used_2),
	.cin(gnd),
	.combout(\ier_wr_en~0_combout ),
	.cout());
defparam \ier_wr_en~0 .lut_mask = 16'hFEFF;
defparam \ier_wr_en~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \always1~0 (
	.dataa(address_2),
	.datab(writedata_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\always1~0_combout ),
	.cout());
defparam \always1~0 .lut_mask = 16'hEEEE;
defparam \always1~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \s_eop~0 (
	.dataa(\set_eop~combout ),
	.datab(\s_eop~q ),
	.datac(\ier_wr_en~0_combout ),
	.datad(\always1~0_combout ),
	.cin(gnd),
	.combout(\s_eop~0_combout ),
	.cout());
defparam \s_eop~0 .lut_mask = 16'hEFFF;
defparam \s_eop~0 .sum_lutc_input = "datac";

dffeas s_eop(
	.clk(clk_clk),
	.d(\s_eop~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\s_eop~q ),
	.prn(vcc));
defparam s_eop.is_wysiwyg = "true";
defparam s_eop.power_up = "low";

fiftyfivenm_lcell_comb \e_eop~0 (
	.dataa(writedata_0),
	.datab(\ier_wr_en~0_combout ),
	.datac(address_2),
	.datad(\e_eop~q ),
	.cin(gnd),
	.combout(\e_eop~0_combout ),
	.cout());
defparam \e_eop~0 .lut_mask = 16'hFF7D;
defparam \e_eop~0 .sum_lutc_input = "datac";

dffeas e_eop(
	.clk(clk_clk),
	.d(\e_eop~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\e_eop~q ),
	.prn(vcc));
defparam e_eop.is_wysiwyg = "true";
defparam e_eop.power_up = "low";

fiftyfivenm_lcell_comb \csr_readdata_nxt[0]~0 (
	.dataa(\s_eop~q ),
	.datab(address_2),
	.datac(gnd),
	.datad(\e_eop~q ),
	.cin(gnd),
	.combout(\csr_readdata_nxt[0]~0_combout ),
	.cout());
defparam \csr_readdata_nxt[0]~0 .lut_mask = 16'h88BB;
defparam \csr_readdata_nxt[0]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \csr_readdata_nxt[0]~2 (
	.dataa(write1),
	.datab(\csr_readdata_nxt[0]~0_combout ),
	.datac(\csr_readdata_nxt[0]~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\csr_readdata_nxt[0]~2_combout ),
	.cout());
defparam \csr_readdata_nxt[0]~2 .lut_mask = 16'hFEFE;
defparam \csr_readdata_nxt[0]~2 .sum_lutc_input = "datac";

dffeas \csr_readdata[0] (
	.clk(clk_clk),
	.d(\csr_readdata_nxt[0]~2_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\csr_readdata[0]~q ),
	.prn(vcc));
defparam \csr_readdata[0] .is_wysiwyg = "true";
defparam \csr_readdata[0] .power_up = "low";

fiftyfivenm_lcell_comb ram_rd_en(
	.dataa(write1),
	.datab(gnd),
	.datac(gnd),
	.datad(address_8),
	.cin(gnd),
	.combout(\ram_rd_en~combout ),
	.cout());
defparam ram_rd_en.lut_mask = 16'hAAFF;
defparam ram_rd_en.sum_lutc_input = "datac";

dffeas ram_rd_en_flp(
	.clk(clk_clk),
	.d(\ram_rd_en~combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ram_rd_en_flp~q ),
	.prn(vcc));
defparam ram_rd_en_flp.is_wysiwyg = "true";
defparam ram_rd_en_flp.power_up = "low";

fiftyfivenm_lcell_comb \readdata_nxt[0]~0 (
	.dataa(\u_ss_ram|altsyncram_component|auto_generated|q_b[0] ),
	.datab(\csr_readdata[0]~q ),
	.datac(gnd),
	.datad(\ram_rd_en_flp~q ),
	.cin(gnd),
	.combout(\readdata_nxt[0]~0_combout ),
	.cout());
defparam \readdata_nxt[0]~0 .lut_mask = 16'hAACC;
defparam \readdata_nxt[0]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \readdata_nxt[2]~1 (
	.dataa(\ram_rd_en_flp~q ),
	.datab(\u_ss_ram|altsyncram_component|auto_generated|q_b[2] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\readdata_nxt[2]~1_combout ),
	.cout());
defparam \readdata_nxt[2]~1 .lut_mask = 16'hEEEE;
defparam \readdata_nxt[2]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \readdata_nxt[1]~2 (
	.dataa(\ram_rd_en_flp~q ),
	.datab(\u_ss_ram|altsyncram_component|auto_generated|q_b[1] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\readdata_nxt[1]~2_combout ),
	.cout());
defparam \readdata_nxt[1]~2 .lut_mask = 16'hEEEE;
defparam \readdata_nxt[1]~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \readdata_nxt[5]~3 (
	.dataa(\ram_rd_en_flp~q ),
	.datab(\u_ss_ram|altsyncram_component|auto_generated|q_b[5] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\readdata_nxt[5]~3_combout ),
	.cout());
defparam \readdata_nxt[5]~3 .lut_mask = 16'hEEEE;
defparam \readdata_nxt[5]~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \readdata_nxt[7]~4 (
	.dataa(\ram_rd_en_flp~q ),
	.datab(\u_ss_ram|altsyncram_component|auto_generated|q_b[7] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\readdata_nxt[7]~4_combout ),
	.cout());
defparam \readdata_nxt[7]~4 .lut_mask = 16'hEEEE;
defparam \readdata_nxt[7]~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \readdata_nxt[6]~5 (
	.dataa(\ram_rd_en_flp~q ),
	.datab(\u_ss_ram|altsyncram_component|auto_generated|q_b[6] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\readdata_nxt[6]~5_combout ),
	.cout());
defparam \readdata_nxt[6]~5 .lut_mask = 16'hEEEE;
defparam \readdata_nxt[6]~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \readdata_nxt[4]~6 (
	.dataa(\ram_rd_en_flp~q ),
	.datab(\u_ss_ram|altsyncram_component|auto_generated|q_b[4] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\readdata_nxt[4]~6_combout ),
	.cout());
defparam \readdata_nxt[4]~6 .lut_mask = 16'hEEEE;
defparam \readdata_nxt[4]~6 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \readdata_nxt[3]~7 (
	.dataa(\ram_rd_en_flp~q ),
	.datab(\u_ss_ram|altsyncram_component|auto_generated|q_b[3] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\readdata_nxt[3]~7_combout ),
	.cout());
defparam \readdata_nxt[3]~7 .lut_mask = 16'hEEEE;
defparam \readdata_nxt[3]~7 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \readdata_nxt[8]~8 (
	.dataa(\ram_rd_en_flp~q ),
	.datab(\u_ss_ram|altsyncram_component|auto_generated|q_b[8] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\readdata_nxt[8]~8_combout ),
	.cout());
defparam \readdata_nxt[8]~8 .lut_mask = 16'hEEEE;
defparam \readdata_nxt[8]~8 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \readdata_nxt[10]~9 (
	.dataa(\ram_rd_en_flp~q ),
	.datab(\u_ss_ram|altsyncram_component|auto_generated|q_b[10] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\readdata_nxt[10]~9_combout ),
	.cout());
defparam \readdata_nxt[10]~9 .lut_mask = 16'hEEEE;
defparam \readdata_nxt[10]~9 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \readdata_nxt[9]~10 (
	.dataa(\ram_rd_en_flp~q ),
	.datab(\u_ss_ram|altsyncram_component|auto_generated|q_b[9] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\readdata_nxt[9]~10_combout ),
	.cout());
defparam \readdata_nxt[9]~10 .lut_mask = 16'hEEEE;
defparam \readdata_nxt[9]~10 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \readdata_nxt[13]~11 (
	.dataa(\ram_rd_en_flp~q ),
	.datab(\u_ss_ram|altsyncram_component|auto_generated|q_b[13] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\readdata_nxt[13]~11_combout ),
	.cout());
defparam \readdata_nxt[13]~11 .lut_mask = 16'hEEEE;
defparam \readdata_nxt[13]~11 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \readdata_nxt[15]~12 (
	.dataa(\ram_rd_en_flp~q ),
	.datab(\u_ss_ram|altsyncram_component|auto_generated|q_b[15] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\readdata_nxt[15]~12_combout ),
	.cout());
defparam \readdata_nxt[15]~12 .lut_mask = 16'hEEEE;
defparam \readdata_nxt[15]~12 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \readdata_nxt[14]~13 (
	.dataa(\ram_rd_en_flp~q ),
	.datab(\u_ss_ram|altsyncram_component|auto_generated|q_b[14] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\readdata_nxt[14]~13_combout ),
	.cout());
defparam \readdata_nxt[14]~13 .lut_mask = 16'hEEEE;
defparam \readdata_nxt[14]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \readdata_nxt[12]~14 (
	.dataa(\ram_rd_en_flp~q ),
	.datab(\u_ss_ram|altsyncram_component|auto_generated|q_b[12] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\readdata_nxt[12]~14_combout ),
	.cout());
defparam \readdata_nxt[12]~14 .lut_mask = 16'hEEEE;
defparam \readdata_nxt[12]~14 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \readdata_nxt[11]~15 (
	.dataa(\ram_rd_en_flp~q ),
	.datab(\u_ss_ram|altsyncram_component|auto_generated|q_b[11] ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\readdata_nxt[11]~15_combout ),
	.cout());
defparam \readdata_nxt[11]~15 .lut_mask = 16'hEEEE;
defparam \readdata_nxt[11]~15 .sum_lutc_input = "datac";

endmodule

module ADC_altera_modular_adc_sample_store_ram (
	q_b_0,
	q_b_2,
	q_b_1,
	q_b_5,
	q_b_7,
	q_b_6,
	q_b_4,
	q_b_3,
	q_b_8,
	slot_num_0,
	slot_num_1,
	slot_num_2,
	slot_num_3,
	slot_num_4,
	slot_num_5,
	q_b_10,
	q_b_9,
	q_b_13,
	q_b_15,
	q_b_14,
	q_b_12,
	q_b_11,
	address_7,
	address_6,
	address_5,
	address_4,
	address_3,
	address_2,
	rsp_valid,
	ram_rd_en,
	rsp_data_0,
	rsp_data_2,
	rsp_data_1,
	rsp_data_5,
	rsp_data_7,
	rsp_data_6,
	rsp_data_4,
	rsp_data_3,
	rsp_data_8,
	rsp_data_10,
	rsp_data_9,
	rsp_data_11,
	GND_port,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_0;
output 	q_b_2;
output 	q_b_1;
output 	q_b_5;
output 	q_b_7;
output 	q_b_6;
output 	q_b_4;
output 	q_b_3;
output 	q_b_8;
input 	slot_num_0;
input 	slot_num_1;
input 	slot_num_2;
input 	slot_num_3;
input 	slot_num_4;
input 	slot_num_5;
output 	q_b_10;
output 	q_b_9;
output 	q_b_13;
output 	q_b_15;
output 	q_b_14;
output 	q_b_12;
output 	q_b_11;
input 	address_7;
input 	address_6;
input 	address_5;
input 	address_4;
input 	address_3;
input 	address_2;
input 	rsp_valid;
input 	ram_rd_en;
input 	rsp_data_0;
input 	rsp_data_2;
input 	rsp_data_1;
input 	rsp_data_5;
input 	rsp_data_7;
input 	rsp_data_6;
input 	rsp_data_4;
input 	rsp_data_3;
input 	rsp_data_8;
input 	rsp_data_10;
input 	rsp_data_9;
input 	rsp_data_11;
input 	GND_port;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ADC_altsyncram_1 altsyncram_component(
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.address_a({slot_num_5,slot_num_4,slot_num_3,slot_num_2,slot_num_1,slot_num_0}),
	.address_b({address_7,address_6,address_5,address_4,address_3,address_2}),
	.wren_a(rsp_valid),
	.rden_b(ram_rd_en),
	.data_a({gnd,gnd,GND_port,gnd,rsp_data_11,rsp_data_10,rsp_data_9,rsp_data_8,rsp_data_7,rsp_data_6,rsp_data_5,rsp_data_4,rsp_data_3,rsp_data_2,rsp_data_1,rsp_data_0}),
	.clock0(clk_clk));

endmodule

module ADC_altsyncram_1 (
	q_b,
	address_a,
	address_b,
	wren_a,
	rden_b,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[5:0] address_a;
input 	[5:0] address_b;
input 	wren_a;
input 	rden_b;
input 	[15:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ADC_altsyncram_v5s1 auto_generated(
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.address_a({address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.wren_a(wren_a),
	.rden_b(rden_b),
	.data_a({data_a[13],data_a[13],data_a[13],data_a[13],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.clock0(clock0));

endmodule

module ADC_altsyncram_v5s1 (
	q_b,
	address_a,
	address_b,
	wren_a,
	rden_b,
	data_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	[5:0] address_a;
input 	[5:0] address_b;
input 	wren_a;
input 	rden_b;
input 	[15:0] data_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

fiftyfivenm_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "ADC_ADC:adc|altera_modular_adc_sample_store:sample_store_internal|altera_modular_adc_sample_store_ram:u_ss_ram|altsyncram:altsyncram_component|altsyncram_v5s1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 6;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 63;
defparam ram_block1a0.port_a_logical_ram_depth = 64;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 6;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 63;
defparam ram_block1a0.port_b_logical_ram_depth = 64;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "ADC_ADC:adc|altera_modular_adc_sample_store:sample_store_internal|altera_modular_adc_sample_store_ram:u_ss_ram|altsyncram:altsyncram_component|altsyncram_v5s1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 6;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 63;
defparam ram_block1a2.port_a_logical_ram_depth = 64;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 6;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 63;
defparam ram_block1a2.port_b_logical_ram_depth = 64;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "ADC_ADC:adc|altera_modular_adc_sample_store:sample_store_internal|altera_modular_adc_sample_store_ram:u_ss_ram|altsyncram:altsyncram_component|altsyncram_v5s1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 6;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 63;
defparam ram_block1a1.port_a_logical_ram_depth = 64;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 6;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 63;
defparam ram_block1a1.port_b_logical_ram_depth = 64;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "ADC_ADC:adc|altera_modular_adc_sample_store:sample_store_internal|altera_modular_adc_sample_store_ram:u_ss_ram|altsyncram:altsyncram_component|altsyncram_v5s1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 6;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 63;
defparam ram_block1a5.port_a_logical_ram_depth = 64;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 6;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 63;
defparam ram_block1a5.port_b_logical_ram_depth = 64;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "ADC_ADC:adc|altera_modular_adc_sample_store:sample_store_internal|altera_modular_adc_sample_store_ram:u_ss_ram|altsyncram:altsyncram_component|altsyncram_v5s1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 6;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 63;
defparam ram_block1a7.port_a_logical_ram_depth = 64;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 6;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 63;
defparam ram_block1a7.port_b_logical_ram_depth = 64;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "ADC_ADC:adc|altera_modular_adc_sample_store:sample_store_internal|altera_modular_adc_sample_store_ram:u_ss_ram|altsyncram:altsyncram_component|altsyncram_v5s1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 6;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 63;
defparam ram_block1a6.port_a_logical_ram_depth = 64;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 6;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 63;
defparam ram_block1a6.port_b_logical_ram_depth = 64;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "ADC_ADC:adc|altera_modular_adc_sample_store:sample_store_internal|altera_modular_adc_sample_store_ram:u_ss_ram|altsyncram:altsyncram_component|altsyncram_v5s1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 6;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 63;
defparam ram_block1a4.port_a_logical_ram_depth = 64;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 6;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 63;
defparam ram_block1a4.port_b_logical_ram_depth = 64;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "ADC_ADC:adc|altera_modular_adc_sample_store:sample_store_internal|altera_modular_adc_sample_store_ram:u_ss_ram|altsyncram:altsyncram_component|altsyncram_v5s1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 6;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 63;
defparam ram_block1a3.port_a_logical_ram_depth = 64;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 6;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 63;
defparam ram_block1a3.port_b_logical_ram_depth = 64;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "ADC_ADC:adc|altera_modular_adc_sample_store:sample_store_internal|altera_modular_adc_sample_store_ram:u_ss_ram|altsyncram:altsyncram_component|altsyncram_v5s1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 6;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 63;
defparam ram_block1a8.port_a_logical_ram_depth = 64;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 6;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 63;
defparam ram_block1a8.port_b_logical_ram_depth = 64;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "ADC_ADC:adc|altera_modular_adc_sample_store:sample_store_internal|altera_modular_adc_sample_store_ram:u_ss_ram|altsyncram:altsyncram_component|altsyncram_v5s1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 6;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 63;
defparam ram_block1a10.port_a_logical_ram_depth = 64;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 6;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 63;
defparam ram_block1a10.port_b_logical_ram_depth = 64;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "ADC_ADC:adc|altera_modular_adc_sample_store:sample_store_internal|altera_modular_adc_sample_store_ram:u_ss_ram|altsyncram:altsyncram_component|altsyncram_v5s1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 6;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 63;
defparam ram_block1a9.port_a_logical_ram_depth = 64;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 6;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 63;
defparam ram_block1a9.port_b_logical_ram_depth = 64;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "ADC_ADC:adc|altera_modular_adc_sample_store:sample_store_internal|altera_modular_adc_sample_store_ram:u_ss_ram|altsyncram:altsyncram_component|altsyncram_v5s1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 6;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 63;
defparam ram_block1a13.port_a_logical_ram_depth = 64;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 6;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 63;
defparam ram_block1a13.port_b_logical_ram_depth = 64;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "ADC_ADC:adc|altera_modular_adc_sample_store:sample_store_internal|altera_modular_adc_sample_store_ram:u_ss_ram|altsyncram:altsyncram_component|altsyncram_v5s1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 6;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 63;
defparam ram_block1a15.port_a_logical_ram_depth = 64;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 6;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 63;
defparam ram_block1a15.port_b_logical_ram_depth = 64;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "ADC_ADC:adc|altera_modular_adc_sample_store:sample_store_internal|altera_modular_adc_sample_store_ram:u_ss_ram|altsyncram:altsyncram_component|altsyncram_v5s1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 6;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 63;
defparam ram_block1a14.port_a_logical_ram_depth = 64;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 6;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 63;
defparam ram_block1a14.port_b_logical_ram_depth = 64;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "ADC_ADC:adc|altera_modular_adc_sample_store:sample_store_internal|altera_modular_adc_sample_store_ram:u_ss_ram|altsyncram:altsyncram_component|altsyncram_v5s1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 6;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 63;
defparam ram_block1a12.port_a_logical_ram_depth = 64;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 6;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 63;
defparam ram_block1a12.port_b_logical_ram_depth = 64;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "M9K";

fiftyfivenm_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "ADC_ADC:adc|altera_modular_adc_sample_store:sample_store_internal|altera_modular_adc_sample_store_ram:u_ss_ram|altsyncram:altsyncram_component|altsyncram_v5s1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 6;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 63;
defparam ram_block1a11.port_a_logical_ram_depth = 64;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 6;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 63;
defparam ram_block1a11.port_b_logical_ram_depth = 64;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "M9K";

endmodule

module ADC_altera_modular_adc_sequencer (
	readdata_0,
	mem_used_1,
	write,
	readdata_2,
	readdata_1,
	readdata_3,
	altera_reset_synchronizer_int_chain_out,
	read,
	src1_valid,
	address_2,
	cmd_ready,
	writedata_0,
	writedata_2,
	writedata_1,
	writedata_3,
	cmd_channel_4,
	cmd_eop,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	readdata_0;
input 	mem_used_1;
input 	write;
output 	readdata_2;
output 	readdata_1;
output 	readdata_3;
input 	altera_reset_synchronizer_int_chain_out;
input 	read;
input 	src1_valid;
input 	address_2;
input 	cmd_ready;
input 	writedata_0;
input 	writedata_2;
input 	writedata_1;
input 	writedata_3;
output 	cmd_channel_4;
output 	cmd_eop;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \u_seq_csr|run~q ;
wire \u_seq_csr|mode[1]~q ;
wire \u_seq_csr|mode[0]~q ;
wire \u_seq_csr|mode[2]~q ;
wire \u_seq_csr|sw_clr_run~q ;
wire \u_seq_ctrl|clr_run~0_combout ;


ADC_altera_modular_adc_sequencer_csr u_seq_csr(
	.readdata_0(readdata_0),
	.mem_used_1(mem_used_1),
	.write(write),
	.readdata_2(readdata_2),
	.readdata_1(readdata_1),
	.readdata_3(readdata_3),
	.rst_n(altera_reset_synchronizer_int_chain_out),
	.read(read),
	.src1_valid(src1_valid),
	.address_2(address_2),
	.run1(\u_seq_csr|run~q ),
	.mode_1(\u_seq_csr|mode[1]~q ),
	.mode_0(\u_seq_csr|mode[0]~q ),
	.mode_2(\u_seq_csr|mode[2]~q ),
	.sw_clr_run1(\u_seq_csr|sw_clr_run~q ),
	.clr_run(\u_seq_ctrl|clr_run~0_combout ),
	.writedata_0(writedata_0),
	.writedata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,writedata_3,writedata_2,writedata_1,gnd}),
	.clk(clk_clk));

ADC_altera_modular_adc_sequencer_ctrl u_seq_ctrl(
	.rst_n(altera_reset_synchronizer_int_chain_out),
	.run(\u_seq_csr|run~q ),
	.mode_1(\u_seq_csr|mode[1]~q ),
	.mode_0(\u_seq_csr|mode[0]~q ),
	.mode_2(\u_seq_csr|mode[2]~q ),
	.sw_clr_run(\u_seq_csr|sw_clr_run~q ),
	.cmd_ready(cmd_ready),
	.clr_run(\u_seq_ctrl|clr_run~0_combout ),
	.cmd_channel_4(cmd_channel_4),
	.cmd_eop1(cmd_eop),
	.clk(clk_clk));

endmodule

module ADC_altera_modular_adc_sequencer_csr (
	readdata_0,
	mem_used_1,
	write,
	readdata_2,
	readdata_1,
	readdata_3,
	rst_n,
	read,
	src1_valid,
	address_2,
	run1,
	mode_1,
	mode_0,
	mode_2,
	sw_clr_run1,
	clr_run,
	writedata_0,
	writedata,
	clk)/* synthesis synthesis_greybox=1 */;
output 	readdata_0;
input 	mem_used_1;
input 	write;
output 	readdata_2;
output 	readdata_1;
output 	readdata_3;
input 	rst_n;
input 	read;
input 	src1_valid;
input 	address_2;
output 	run1;
output 	mode_1;
output 	mode_0;
output 	mode_2;
output 	sw_clr_run1;
input 	clr_run;
input 	writedata_0;
input 	[31:0] writedata;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \cmd_rd_en~0_combout ;
wire \readdata_nxt[0]~combout ;
wire \readdata_nxt[2]~combout ;
wire \readdata_nxt[1]~combout ;
wire \readdata_nxt[3]~combout ;
wire \always0~0_combout ;
wire \run~0_combout ;
wire \always0~1_combout ;
wire \Equal1~0_combout ;
wire \sw_clr_run~0_combout ;
wire \sw_clr_run~1_combout ;


dffeas \readdata[0] (
	.clk(clk),
	.d(\readdata_nxt[0]~combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk),
	.d(\readdata_nxt[2]~combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk),
	.d(\readdata_nxt[1]~combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[3] (
	.clk(clk),
	.d(\readdata_nxt[3]~combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas run(
	.clk(clk),
	.d(\run~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(run1),
	.prn(vcc));
defparam run.is_wysiwyg = "true";
defparam run.power_up = "low";

dffeas \mode[1] (
	.clk(clk),
	.d(writedata[2]),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(mode_1),
	.prn(vcc));
defparam \mode[1] .is_wysiwyg = "true";
defparam \mode[1] .power_up = "low";

dffeas \mode[0] (
	.clk(clk),
	.d(writedata[1]),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(mode_0),
	.prn(vcc));
defparam \mode[0] .is_wysiwyg = "true";
defparam \mode[0] .power_up = "low";

dffeas \mode[2] (
	.clk(clk),
	.d(writedata[3]),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~1_combout ),
	.q(mode_2),
	.prn(vcc));
defparam \mode[2] .is_wysiwyg = "true";
defparam \mode[2] .power_up = "low";

dffeas sw_clr_run(
	.clk(clk),
	.d(\sw_clr_run~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sw_clr_run1),
	.prn(vcc));
defparam sw_clr_run.is_wysiwyg = "true";
defparam sw_clr_run.power_up = "low";

fiftyfivenm_lcell_comb \cmd_rd_en~0 (
	.dataa(write),
	.datab(read),
	.datac(mem_used_1),
	.datad(address_2),
	.cin(gnd),
	.combout(\cmd_rd_en~0_combout ),
	.cout());
defparam \cmd_rd_en~0 .lut_mask = 16'hEFFF;
defparam \cmd_rd_en~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \readdata_nxt[0] (
	.dataa(read),
	.datab(src1_valid),
	.datac(\cmd_rd_en~0_combout ),
	.datad(run1),
	.cin(gnd),
	.combout(\readdata_nxt[0]~combout ),
	.cout());
defparam \readdata_nxt[0] .lut_mask = 16'hFFFE;
defparam \readdata_nxt[0] .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \readdata_nxt[2] (
	.dataa(read),
	.datab(src1_valid),
	.datac(\cmd_rd_en~0_combout ),
	.datad(mode_1),
	.cin(gnd),
	.combout(\readdata_nxt[2]~combout ),
	.cout());
defparam \readdata_nxt[2] .lut_mask = 16'hFFFE;
defparam \readdata_nxt[2] .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \readdata_nxt[1] (
	.dataa(read),
	.datab(src1_valid),
	.datac(\cmd_rd_en~0_combout ),
	.datad(mode_0),
	.cin(gnd),
	.combout(\readdata_nxt[1]~combout ),
	.cout());
defparam \readdata_nxt[1] .lut_mask = 16'hFFFE;
defparam \readdata_nxt[1] .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \readdata_nxt[3] (
	.dataa(read),
	.datab(src1_valid),
	.datac(\cmd_rd_en~0_combout ),
	.datad(mode_2),
	.cin(gnd),
	.combout(\readdata_nxt[3]~combout ),
	.cout());
defparam \readdata_nxt[3] .lut_mask = 16'hFFFE;
defparam \readdata_nxt[3] .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \always0~0 (
	.dataa(write),
	.datab(src1_valid),
	.datac(\cmd_rd_en~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
defparam \always0~0 .lut_mask = 16'hFEFE;
defparam \always0~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \run~0 (
	.dataa(clr_run),
	.datab(run1),
	.datac(writedata_0),
	.datad(\always0~0_combout ),
	.cin(gnd),
	.combout(\run~0_combout ),
	.cout());
defparam \run~0 .lut_mask = 16'hFFFE;
defparam \run~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \always0~1 (
	.dataa(write),
	.datab(src1_valid),
	.datac(\cmd_rd_en~0_combout ),
	.datad(run1),
	.cin(gnd),
	.combout(\always0~1_combout ),
	.cout());
defparam \always0~1 .lut_mask = 16'hFEFF;
defparam \always0~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Equal1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(mode_1),
	.datad(mode_2),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
defparam \Equal1~0 .lut_mask = 16'h0FFF;
defparam \Equal1~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \sw_clr_run~0 (
	.dataa(run1),
	.datab(\Equal1~0_combout ),
	.datac(mode_0),
	.datad(writedata_0),
	.cin(gnd),
	.combout(\sw_clr_run~0_combout ),
	.cout());
defparam \sw_clr_run~0 .lut_mask = 16'hEFFF;
defparam \sw_clr_run~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \sw_clr_run~1 (
	.dataa(clr_run),
	.datab(sw_clr_run1),
	.datac(\always0~0_combout ),
	.datad(\sw_clr_run~0_combout ),
	.cin(gnd),
	.combout(\sw_clr_run~1_combout ),
	.cout());
defparam \sw_clr_run~1 .lut_mask = 16'hFFFE;
defparam \sw_clr_run~1 .sum_lutc_input = "datac";

endmodule

module ADC_altera_modular_adc_sequencer_ctrl (
	rst_n,
	run,
	mode_1,
	mode_0,
	mode_2,
	sw_clr_run,
	cmd_ready,
	clr_run,
	cmd_channel_4,
	cmd_eop1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	rst_n;
input 	run;
input 	mode_1;
input 	mode_0;
input 	mode_2;
input 	sw_clr_run;
input 	cmd_ready;
output 	clr_run;
output 	cmd_channel_4;
output 	cmd_eop1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \valid_req~0_combout ;
wire \cmd_eop~0_combout ;
wire \cmd_eop~1_combout ;
wire \seq_state_nxt~0_combout ;
wire \seq_state~q ;
wire \valid_req~1_combout ;
wire \cmd_channel~0_combout ;
wire \cmd_eop~2_combout ;


fiftyfivenm_lcell_comb \clr_run~0 (
	.dataa(\valid_req~0_combout ),
	.datab(gnd),
	.datac(cmd_ready),
	.datad(\seq_state~q ),
	.cin(gnd),
	.combout(clr_run),
	.cout());
defparam \clr_run~0 .lut_mask = 16'hAFFF;
defparam \clr_run~0 .sum_lutc_input = "datac";

dffeas \cmd_channel[4] (
	.clk(clk),
	.d(\cmd_channel~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\cmd_eop~2_combout ),
	.q(cmd_channel_4),
	.prn(vcc));
defparam \cmd_channel[4] .is_wysiwyg = "true";
defparam \cmd_channel[4] .power_up = "low";

dffeas cmd_eop(
	.clk(clk),
	.d(\valid_req~1_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\cmd_eop~2_combout ),
	.q(cmd_eop1),
	.prn(vcc));
defparam cmd_eop.is_wysiwyg = "true";
defparam cmd_eop.power_up = "low";

fiftyfivenm_lcell_comb \valid_req~0 (
	.dataa(mode_1),
	.datab(mode_2),
	.datac(mode_0),
	.datad(sw_clr_run),
	.cin(gnd),
	.combout(\valid_req~0_combout ),
	.cout());
defparam \valid_req~0 .lut_mask = 16'h6FFF;
defparam \valid_req~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \cmd_eop~0 (
	.dataa(mode_0),
	.datab(mode_1),
	.datac(mode_2),
	.datad(gnd),
	.cin(gnd),
	.combout(\cmd_eop~0_combout ),
	.cout());
defparam \cmd_eop~0 .lut_mask = 16'hBEBE;
defparam \cmd_eop~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \cmd_eop~1 (
	.dataa(run),
	.datab(\cmd_eop~0_combout ),
	.datac(gnd),
	.datad(\seq_state~q ),
	.cin(gnd),
	.combout(\cmd_eop~1_combout ),
	.cout());
defparam \cmd_eop~1 .lut_mask = 16'hEEFF;
defparam \cmd_eop~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \seq_state_nxt~0 (
	.dataa(\cmd_eop~1_combout ),
	.datab(\seq_state~q ),
	.datac(\valid_req~0_combout ),
	.datad(cmd_ready),
	.cin(gnd),
	.combout(\seq_state_nxt~0_combout ),
	.cout());
defparam \seq_state_nxt~0 .lut_mask = 16'hFEFF;
defparam \seq_state_nxt~0 .sum_lutc_input = "datac";

dffeas seq_state(
	.clk(clk),
	.d(\seq_state_nxt~0_combout ),
	.asdata(vcc),
	.clrn(rst_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\seq_state~q ),
	.prn(vcc));
defparam seq_state.is_wysiwyg = "true";
defparam seq_state.power_up = "low";

fiftyfivenm_lcell_comb \valid_req~1 (
	.dataa(\cmd_eop~1_combout ),
	.datab(\valid_req~0_combout ),
	.datac(cmd_ready),
	.datad(\seq_state~q ),
	.cin(gnd),
	.combout(\valid_req~1_combout ),
	.cout());
defparam \valid_req~1 .lut_mask = 16'hFFFE;
defparam \valid_req~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \cmd_channel~0 (
	.dataa(mode_1),
	.datab(mode_0),
	.datac(mode_2),
	.datad(\valid_req~1_combout ),
	.cin(gnd),
	.combout(\cmd_channel~0_combout ),
	.cout());
defparam \cmd_channel~0 .lut_mask = 16'hFFFE;
defparam \cmd_channel~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \cmd_eop~2 (
	.dataa(cmd_ready),
	.datab(run),
	.datac(\cmd_eop~0_combout ),
	.datad(\seq_state~q ),
	.cin(gnd),
	.combout(\cmd_eop~2_combout ),
	.cout());
defparam \cmd_eop~2 .lut_mask = 16'hFEFF;
defparam \cmd_eop~2 .sum_lutc_input = "datac";

endmodule

module ADC_ADC_AvalonBridge (
	tdo,
	read_latency_shift_reg_1,
	src_data_0,
	address_7,
	address_6,
	address_5,
	address_4,
	address_9,
	address_3,
	address_8,
	master_write,
	av_waitrequest,
	src_data_2,
	src_data_1,
	src_payload,
	readdata_7,
	src_payload1,
	src_payload2,
	src_data_3,
	src_payload3,
	master_read,
	address_2,
	WideOr1,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	writedata_0,
	writedata_2,
	writedata_1,
	writedata_3,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	splitter_nodes_receive_0_3,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	irf_reg_0_1,
	irf_reg_1_1,
	irf_reg_2_1,
	clk_clk,
	reset_reset_n)/* synthesis synthesis_greybox=1 */;
output 	tdo;
input 	read_latency_shift_reg_1;
input 	src_data_0;
output 	address_7;
output 	address_6;
output 	address_5;
output 	address_4;
output 	address_9;
output 	address_3;
output 	address_8;
output 	master_write;
input 	av_waitrequest;
input 	src_data_2;
input 	src_data_1;
input 	src_payload;
input 	readdata_7;
input 	src_payload1;
input 	src_payload2;
input 	src_data_3;
input 	src_payload3;
output 	master_read;
output 	address_2;
input 	WideOr1;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
output 	writedata_0;
output 	writedata_2;
output 	writedata_1;
output 	writedata_3;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	splitter_nodes_receive_0_3;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	clk_clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \transacto|p2m|out_endofpacket~q ;
wire \rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \p2b|out_data[0]~q ;
wire \p2b|out_valid~q ;
wire \jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|sink_crosser|in_data_toggle~q ;
wire \jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|sink_crosser|out_to_in_synchronizer|dreg[6]~q ;
wire \p2b|out_data[2]~q ;
wire \p2b|out_data[1]~q ;
wire \p2b|out_data[6]~q ;
wire \p2b|out_data[7]~q ;
wire \p2b|out_data[5]~q ;
wire \p2b|out_data[3]~q ;
wire \p2b|out_data[4]~q ;
wire \transacto|p2m|out_data[0]~q ;
wire \transacto|p2m|out_startofpacket~q ;
wire \transacto|p2m|out_data[2]~q ;
wire \transacto|p2m|out_data[1]~q ;
wire \transacto|p2m|out_data[5]~q ;
wire \transacto|p2m|out_data[7]~q ;
wire \transacto|p2m|out_data[6]~q ;
wire \transacto|p2m|out_data[4]~q ;
wire \transacto|p2m|out_data[3]~q ;
wire \transacto|p2m|out_valid~q ;
wire \b2p|received_esc~q ;
wire \fifo|out_payload[3]~q ;
wire \fifo|out_payload[6]~q ;
wire \fifo|out_payload[5]~q ;
wire \fifo|out_payload[4]~q ;
wire \fifo|out_payload[7]~q ;
wire \fifo|out_payload[1]~q ;
wire \fifo|out_payload[2]~q ;
wire \b2p|out_valid~0_combout ;
wire \fifo|out_valid~q ;
wire \transacto|p2m|in_ready_0~q ;
wire \transacto|p2m|enable~0_combout ;
wire \b2p|out_channel[0]~q ;
wire \b2p|out_channel[7]~q ;
wire \b2p|out_channel[6]~q ;
wire \b2p|out_channel[5]~q ;
wire \b2p|out_channel[4]~q ;
wire \b2p|out_channel[3]~q ;
wire \b2p|out_channel[2]~q ;
wire \b2p|out_channel[1]~q ;
wire \b2p|received_channel~q ;
wire \p2b|in_ready~combout ;
wire \b2p|out_startofpacket~q ;
wire \b2p|out_endofpacket~q ;
wire \fifo|out_payload[0]~q ;
wire \b2p|out_data[5]~0_combout ;
wire \jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|source_crosser|src_valid~q ;
wire \jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|source_crosser|src_data[3]~q ;
wire \jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|source_crosser|src_data[6]~q ;
wire \jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|source_crosser|src_data[5]~q ;
wire \jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|source_crosser|src_data[4]~q ;
wire \jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|source_crosser|src_data[7]~q ;
wire \jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|source_crosser|src_data[1]~q ;
wire \jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|source_crosser|src_data[2]~q ;
wire \jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|source_crosser|src_data[0]~q ;


ADC_altera_avalon_packets_to_master transacto(
	.out_endofpacket(\transacto|p2m|out_endofpacket~q ),
	.altera_reset_synchronizer_int_chain_out(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.out_data_0(\transacto|p2m|out_data[0]~q ),
	.out_startofpacket(\transacto|p2m|out_startofpacket~q ),
	.out_data_2(\transacto|p2m|out_data[2]~q ),
	.out_data_1(\transacto|p2m|out_data[1]~q ),
	.out_data_5(\transacto|p2m|out_data[5]~q ),
	.out_data_7(\transacto|p2m|out_data[7]~q ),
	.out_data_6(\transacto|p2m|out_data[6]~q ),
	.out_data_4(\transacto|p2m|out_data[4]~q ),
	.out_data_3(\transacto|p2m|out_data[3]~q ),
	.out_valid(\transacto|p2m|out_valid~q ),
	.read_latency_shift_reg_1(read_latency_shift_reg_1),
	.src_data_0(src_data_0),
	.address_7(address_7),
	.address_6(address_6),
	.address_5(address_5),
	.address_4(address_4),
	.address_9(address_9),
	.address_3(address_3),
	.address_8(address_8),
	.write(master_write),
	.av_waitrequest(av_waitrequest),
	.received_esc(\b2p|received_esc~q ),
	.out_payload_3(\fifo|out_payload[3]~q ),
	.out_payload_6(\fifo|out_payload[6]~q ),
	.out_payload_5(\fifo|out_payload[5]~q ),
	.out_payload_4(\fifo|out_payload[4]~q ),
	.out_payload_7(\fifo|out_payload[7]~q ),
	.out_payload_1(\fifo|out_payload[1]~q ),
	.out_payload_2(\fifo|out_payload[2]~q ),
	.out_valid1(\b2p|out_valid~0_combout ),
	.out_valid2(\fifo|out_valid~q ),
	.in_ready_0(\transacto|p2m|in_ready_0~q ),
	.enable(\transacto|p2m|enable~0_combout ),
	.out_channel_0(\b2p|out_channel[0]~q ),
	.out_channel_7(\b2p|out_channel[7]~q ),
	.out_channel_6(\b2p|out_channel[6]~q ),
	.out_channel_5(\b2p|out_channel[5]~q ),
	.out_channel_4(\b2p|out_channel[4]~q ),
	.out_channel_3(\b2p|out_channel[3]~q ),
	.out_channel_2(\b2p|out_channel[2]~q ),
	.out_channel_1(\b2p|out_channel[1]~q ),
	.received_channel(\b2p|received_channel~q ),
	.in_ready(\p2b|in_ready~combout ),
	.src_data_2(src_data_2),
	.src_data_1(src_data_1),
	.src_payload(src_payload),
	.readdata_7(readdata_7),
	.src_payload1(src_payload1),
	.src_payload2(src_payload2),
	.src_data_3(src_data_3),
	.src_payload3(src_payload3),
	.read(master_read),
	.address_2(address_2),
	.WideOr1(WideOr1),
	.out_startofpacket1(\b2p|out_startofpacket~q ),
	.out_endofpacket1(\b2p|out_endofpacket~q ),
	.out_payload_0(\fifo|out_payload[0]~q ),
	.out_data_51(\b2p|out_data[5]~0_combout ),
	.src_payload4(src_payload4),
	.src_payload5(src_payload5),
	.src_payload6(src_payload6),
	.src_payload7(src_payload7),
	.src_payload8(src_payload8),
	.src_payload9(src_payload9),
	.src_payload10(src_payload10),
	.writedata_0(writedata_0),
	.writedata_2(writedata_2),
	.writedata_1(writedata_1),
	.writedata_3(writedata_3),
	.clk_clk(clk_clk));

ADC_altera_avalon_st_packets_to_bytes p2b(
	.out_endofpacket(\transacto|p2m|out_endofpacket~q ),
	.reset_n(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.out_data_0(\p2b|out_data[0]~q ),
	.out_valid1(\p2b|out_valid~q ),
	.in_data_toggle(\jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|sink_crosser|in_data_toggle~q ),
	.dreg_6(\jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|sink_crosser|out_to_in_synchronizer|dreg[6]~q ),
	.out_data_2(\p2b|out_data[2]~q ),
	.out_data_1(\p2b|out_data[1]~q ),
	.out_data_6(\p2b|out_data[6]~q ),
	.out_data_7(\p2b|out_data[7]~q ),
	.out_data_5(\p2b|out_data[5]~q ),
	.out_data_3(\p2b|out_data[3]~q ),
	.out_data_4(\p2b|out_data[4]~q ),
	.out_data_01(\transacto|p2m|out_data[0]~q ),
	.out_startofpacket(\transacto|p2m|out_startofpacket~q ),
	.out_data_21(\transacto|p2m|out_data[2]~q ),
	.out_data_11(\transacto|p2m|out_data[1]~q ),
	.out_data_51(\transacto|p2m|out_data[5]~q ),
	.out_data_71(\transacto|p2m|out_data[7]~q ),
	.out_data_61(\transacto|p2m|out_data[6]~q ),
	.out_data_41(\transacto|p2m|out_data[4]~q ),
	.out_data_31(\transacto|p2m|out_data[3]~q ),
	.out_valid2(\transacto|p2m|out_valid~q ),
	.in_ready1(\p2b|in_ready~combout ),
	.clk(clk_clk));

ADC_altera_avalon_st_bytes_to_packets b2p(
	.reset_n(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.received_esc1(\b2p|received_esc~q ),
	.out_payload_3(\fifo|out_payload[3]~q ),
	.out_payload_6(\fifo|out_payload[6]~q ),
	.out_payload_5(\fifo|out_payload[5]~q ),
	.out_payload_4(\fifo|out_payload[4]~q ),
	.out_payload_7(\fifo|out_payload[7]~q ),
	.out_payload_1(\fifo|out_payload[1]~q ),
	.out_payload_2(\fifo|out_payload[2]~q ),
	.out_valid(\b2p|out_valid~0_combout ),
	.out_valid1(\fifo|out_valid~q ),
	.in_ready_0(\transacto|p2m|in_ready_0~q ),
	.enable(\transacto|p2m|enable~0_combout ),
	.out_channel_0(\b2p|out_channel[0]~q ),
	.out_channel_7(\b2p|out_channel[7]~q ),
	.out_channel_6(\b2p|out_channel[6]~q ),
	.out_channel_5(\b2p|out_channel[5]~q ),
	.out_channel_4(\b2p|out_channel[4]~q ),
	.out_channel_3(\b2p|out_channel[3]~q ),
	.out_channel_2(\b2p|out_channel[2]~q ),
	.out_channel_1(\b2p|out_channel[1]~q ),
	.received_channel1(\b2p|received_channel~q ),
	.out_startofpacket1(\b2p|out_startofpacket~q ),
	.out_endofpacket1(\b2p|out_endofpacket~q ),
	.out_payload_0(\fifo|out_payload[0]~q ),
	.out_data_5(\b2p|out_data[5]~0_combout ),
	.clk(clk_clk));

ADC_altera_avalon_sc_fifo fifo(
	.reset(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.out_payload_3(\fifo|out_payload[3]~q ),
	.out_payload_6(\fifo|out_payload[6]~q ),
	.out_payload_5(\fifo|out_payload[5]~q ),
	.out_payload_4(\fifo|out_payload[4]~q ),
	.out_payload_7(\fifo|out_payload[7]~q ),
	.out_payload_1(\fifo|out_payload[1]~q ),
	.out_payload_2(\fifo|out_payload[2]~q ),
	.out_valid1(\fifo|out_valid~q ),
	.in_ready_0(\transacto|p2m|in_ready_0~q ),
	.out_payload_0(\fifo|out_payload[0]~q ),
	.src_valid(\jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|source_crosser|src_valid~q ),
	.src_data_3(\jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|source_crosser|src_data[3]~q ),
	.src_data_6(\jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|source_crosser|src_data[6]~q ),
	.src_data_5(\jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|source_crosser|src_data[5]~q ),
	.src_data_4(\jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|source_crosser|src_data[4]~q ),
	.src_data_7(\jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|source_crosser|src_data[7]~q ),
	.src_data_1(\jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|source_crosser|src_data[1]~q ),
	.src_data_2(\jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|source_crosser|src_data[2]~q ),
	.src_data_0(\jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|source_crosser|src_data[0]~q ),
	.clk(clk_clk));

ADC_altera_reset_controller rst_controller(
	.altera_reset_synchronizer_int_chain_out(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.clk_clk(clk_clk),
	.reset_reset_n(reset_reset_n));

ADC_altera_avalon_st_jtag_interface jtag_phy_embedded_in_jtag_master(
	.tdo(tdo),
	.altera_reset_synchronizer_int_chain_out(\rst_controller|alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.out_data_0(\p2b|out_data[0]~q ),
	.out_valid(\p2b|out_valid~q ),
	.in_data_toggle(\jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|sink_crosser|in_data_toggle~q ),
	.dreg_6(\jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|sink_crosser|out_to_in_synchronizer|dreg[6]~q ),
	.out_data_2(\p2b|out_data[2]~q ),
	.out_data_1(\p2b|out_data[1]~q ),
	.out_data_6(\p2b|out_data[6]~q ),
	.out_data_7(\p2b|out_data[7]~q ),
	.out_data_5(\p2b|out_data[5]~q ),
	.out_data_3(\p2b|out_data[3]~q ),
	.out_data_4(\p2b|out_data[4]~q ),
	.src_valid(\jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|source_crosser|src_valid~q ),
	.src_data_3(\jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|source_crosser|src_data[3]~q ),
	.src_data_6(\jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|source_crosser|src_data[6]~q ),
	.src_data_5(\jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|source_crosser|src_data[5]~q ),
	.src_data_4(\jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|source_crosser|src_data[4]~q ),
	.src_data_7(\jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|source_crosser|src_data[7]~q ),
	.src_data_1(\jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|source_crosser|src_data[1]~q ),
	.src_data_2(\jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|source_crosser|src_data[2]~q ),
	.src_data_0(\jtag_phy_embedded_in_jtag_master|normal.jtag_dc_streaming|source_crosser|src_data[0]~q ),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.splitter_nodes_receive_0_3(splitter_nodes_receive_0_3),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.irf_reg_0_1(irf_reg_0_1),
	.irf_reg_1_1(irf_reg_1_1),
	.irf_reg_2_1(irf_reg_2_1),
	.clk_clk(clk_clk));

endmodule

module ADC_altera_avalon_packets_to_master (
	out_endofpacket,
	altera_reset_synchronizer_int_chain_out,
	out_data_0,
	out_startofpacket,
	out_data_2,
	out_data_1,
	out_data_5,
	out_data_7,
	out_data_6,
	out_data_4,
	out_data_3,
	out_valid,
	read_latency_shift_reg_1,
	src_data_0,
	address_7,
	address_6,
	address_5,
	address_4,
	address_9,
	address_3,
	address_8,
	write,
	av_waitrequest,
	received_esc,
	out_payload_3,
	out_payload_6,
	out_payload_5,
	out_payload_4,
	out_payload_7,
	out_payload_1,
	out_payload_2,
	out_valid1,
	out_valid2,
	in_ready_0,
	enable,
	out_channel_0,
	out_channel_7,
	out_channel_6,
	out_channel_5,
	out_channel_4,
	out_channel_3,
	out_channel_2,
	out_channel_1,
	received_channel,
	in_ready,
	src_data_2,
	src_data_1,
	src_payload,
	readdata_7,
	src_payload1,
	src_payload2,
	src_data_3,
	src_payload3,
	read,
	address_2,
	WideOr1,
	out_startofpacket1,
	out_endofpacket1,
	out_payload_0,
	out_data_51,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	writedata_0,
	writedata_2,
	writedata_1,
	writedata_3,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	out_endofpacket;
input 	altera_reset_synchronizer_int_chain_out;
output 	out_data_0;
output 	out_startofpacket;
output 	out_data_2;
output 	out_data_1;
output 	out_data_5;
output 	out_data_7;
output 	out_data_6;
output 	out_data_4;
output 	out_data_3;
output 	out_valid;
input 	read_latency_shift_reg_1;
input 	src_data_0;
output 	address_7;
output 	address_6;
output 	address_5;
output 	address_4;
output 	address_9;
output 	address_3;
output 	address_8;
output 	write;
input 	av_waitrequest;
input 	received_esc;
input 	out_payload_3;
input 	out_payload_6;
input 	out_payload_5;
input 	out_payload_4;
input 	out_payload_7;
input 	out_payload_1;
input 	out_payload_2;
input 	out_valid1;
input 	out_valid2;
output 	in_ready_0;
output 	enable;
input 	out_channel_0;
input 	out_channel_7;
input 	out_channel_6;
input 	out_channel_5;
input 	out_channel_4;
input 	out_channel_3;
input 	out_channel_2;
input 	out_channel_1;
input 	received_channel;
input 	in_ready;
input 	src_data_2;
input 	src_data_1;
input 	src_payload;
input 	readdata_7;
input 	src_payload1;
input 	src_payload2;
input 	src_data_3;
input 	src_payload3;
output 	read;
output 	address_2;
input 	WideOr1;
input 	out_startofpacket1;
input 	out_endofpacket1;
input 	out_payload_0;
input 	out_data_51;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
output 	writedata_0;
output 	writedata_2;
output 	writedata_1;
output 	writedata_3;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ADC_packets_to_master p2m(
	.out_endofpacket1(out_endofpacket),
	.reset_n(altera_reset_synchronizer_int_chain_out),
	.out_data_0(out_data_0),
	.out_startofpacket1(out_startofpacket),
	.out_data_2(out_data_2),
	.out_data_1(out_data_1),
	.out_data_5(out_data_5),
	.out_data_7(out_data_7),
	.out_data_6(out_data_6),
	.out_data_4(out_data_4),
	.out_data_3(out_data_3),
	.out_valid1(out_valid),
	.read_latency_shift_reg_1(read_latency_shift_reg_1),
	.src_data_0(src_data_0),
	.address_7(address_7),
	.address_6(address_6),
	.address_5(address_5),
	.address_4(address_4),
	.address_9(address_9),
	.address_3(address_3),
	.address_8(address_8),
	.write1(write),
	.av_waitrequest(av_waitrequest),
	.received_esc(received_esc),
	.in_data({out_payload_7,out_payload_6,out_data_51,out_payload_4,out_payload_3,out_payload_2,out_payload_1,out_payload_0}),
	.out_payload_5(out_payload_5),
	.out_valid2(out_valid1),
	.out_valid3(out_valid2),
	.in_ready_01(in_ready_0),
	.enable1(enable),
	.out_channel_0(out_channel_0),
	.out_channel_7(out_channel_7),
	.out_channel_6(out_channel_6),
	.out_channel_5(out_channel_5),
	.out_channel_4(out_channel_4),
	.out_channel_3(out_channel_3),
	.out_channel_2(out_channel_2),
	.out_channel_1(out_channel_1),
	.received_channel(received_channel),
	.in_ready(in_ready),
	.src_data_2(src_data_2),
	.src_data_1(src_data_1),
	.src_payload(src_payload),
	.readdata_7(readdata_7),
	.src_payload1(src_payload1),
	.src_payload2(src_payload2),
	.src_data_3(src_data_3),
	.readdata({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_payload7,src_payload8,src_payload6,src_payload9,src_payload10,src_payload4,src_payload5,src_payload3,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.read1(read),
	.address_2(address_2),
	.WideOr1(WideOr1),
	.out_startofpacket2(out_startofpacket1),
	.out_endofpacket2(out_endofpacket1),
	.writedata_0(writedata_0),
	.writedata_2(writedata_2),
	.writedata_1(writedata_1),
	.writedata_3(writedata_3),
	.clk(clk_clk));

endmodule

module ADC_packets_to_master (
	out_endofpacket1,
	reset_n,
	out_data_0,
	out_startofpacket1,
	out_data_2,
	out_data_1,
	out_data_5,
	out_data_7,
	out_data_6,
	out_data_4,
	out_data_3,
	out_valid1,
	read_latency_shift_reg_1,
	src_data_0,
	address_7,
	address_6,
	address_5,
	address_4,
	address_9,
	address_3,
	address_8,
	write1,
	av_waitrequest,
	received_esc,
	in_data,
	out_payload_5,
	out_valid2,
	out_valid3,
	in_ready_01,
	enable1,
	out_channel_0,
	out_channel_7,
	out_channel_6,
	out_channel_5,
	out_channel_4,
	out_channel_3,
	out_channel_2,
	out_channel_1,
	received_channel,
	in_ready,
	src_data_2,
	src_data_1,
	src_payload,
	readdata_7,
	src_payload1,
	src_payload2,
	src_data_3,
	readdata,
	read1,
	address_2,
	WideOr1,
	out_startofpacket2,
	out_endofpacket2,
	writedata_0,
	writedata_2,
	writedata_1,
	writedata_3,
	clk)/* synthesis synthesis_greybox=1 */;
output 	out_endofpacket1;
input 	reset_n;
output 	out_data_0;
output 	out_startofpacket1;
output 	out_data_2;
output 	out_data_1;
output 	out_data_5;
output 	out_data_7;
output 	out_data_6;
output 	out_data_4;
output 	out_data_3;
output 	out_valid1;
input 	read_latency_shift_reg_1;
input 	src_data_0;
output 	address_7;
output 	address_6;
output 	address_5;
output 	address_4;
output 	address_9;
output 	address_3;
output 	address_8;
output 	write1;
input 	av_waitrequest;
input 	received_esc;
input 	[7:0] in_data;
input 	out_payload_5;
input 	out_valid2;
input 	out_valid3;
output 	in_ready_01;
output 	enable1;
input 	out_channel_0;
input 	out_channel_7;
input 	out_channel_6;
input 	out_channel_5;
input 	out_channel_4;
input 	out_channel_3;
input 	out_channel_2;
input 	out_channel_1;
input 	received_channel;
input 	in_ready;
input 	src_data_2;
input 	src_data_1;
input 	src_payload;
input 	readdata_7;
input 	src_payload1;
input 	src_payload2;
input 	src_data_3;
input 	[31:0] readdata;
output 	read1;
output 	address_2;
input 	WideOr1;
input 	out_startofpacket2;
input 	out_endofpacket2;
output 	writedata_0;
output 	writedata_2;
output 	writedata_1;
output 	writedata_3;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \enable~1_combout ;
wire \enable~2_combout ;
wire \enable~3_combout ;
wire \enable~combout ;
wire \always1~0_combout ;
wire \command[7]~q ;
wire \command[6]~q ;
wire \command[5]~q ;
wire \command[3]~q ;
wire \Equal2~0_combout ;
wire \command[0]~q ;
wire \command[1]~q ;
wire \Equal2~1_combout ;
wire \Selector72~1_combout ;
wire \Selector39~0_combout ;
wire \last_trans~q ;
wire \state~59_combout ;
wire \state~79_combout ;
wire \state~60_combout ;
wire \state.RETURN_PACKET~q ;
wire \Add0~0_combout ;
wire \command[4]~q ;
wire \counter~16_combout ;
wire \counter[0]~15_combout ;
wire \Add3~0_combout ;
wire \out_data[0]~7_combout ;
wire \state~61_combout ;
wire \address[9]~2_combout ;
wire \state~71_combout ;
wire \state~80_combout ;
wire \state.READ_ASSERT~q ;
wire \state~49_combout ;
wire \state~58_combout ;
wire \state~78_combout ;
wire \state.READ_DATA_WAIT~q ;
wire \current_byte[1]~0_combout ;
wire \state~50_combout ;
wire \state~51_combout ;
wire \state~52_combout ;
wire \state~53_combout ;
wire \write~0_combout ;
wire \in_ready_0~0_combout ;
wire \in_ready_0~1_combout ;
wire \state~54_combout ;
wire \state~55_combout ;
wire \state~56_combout ;
wire \state~57_combout ;
wire \state.READ_CMD_WAIT~q ;
wire \out_data~4_combout ;
wire \state~62_combout ;
wire \state.READ_SEND_ISSUE~q ;
wire \state~70_combout ;
wire \state.READ_SEND_WAIT~q ;
wire \counter[9]~17_combout ;
wire \counter[4]~19_combout ;
wire \counter[0]~q ;
wire \Add0~1 ;
wire \Add0~2_combout ;
wire \counter~26_combout ;
wire \counter[1]~14_combout ;
wire \Add3~1 ;
wire \Add3~2_combout ;
wire \counter[1]~q ;
wire \Add0~3 ;
wire \Add0~4_combout ;
wire \counter~25_combout ;
wire \counter[2]~13_combout ;
wire \Add3~3 ;
wire \Add3~4_combout ;
wire \counter[2]~q ;
wire \Add0~5 ;
wire \Add0~6_combout ;
wire \counter~24_combout ;
wire \counter[3]~12_combout ;
wire \Add3~5 ;
wire \Add3~6_combout ;
wire \counter[3]~q ;
wire \Add0~7 ;
wire \Add0~8_combout ;
wire \counter~23_combout ;
wire \counter[4]~11_combout ;
wire \Add3~7 ;
wire \Add3~8_combout ;
wire \counter[4]~q ;
wire \Add0~9 ;
wire \Add0~10_combout ;
wire \counter~22_combout ;
wire \counter[5]~10_combout ;
wire \Add3~9 ;
wire \Add3~10_combout ;
wire \counter[5]~q ;
wire \Add0~11 ;
wire \Add0~12_combout ;
wire \counter~21_combout ;
wire \counter[6]~9_combout ;
wire \Add3~11 ;
wire \Add3~12_combout ;
wire \counter[6]~q ;
wire \Add0~13 ;
wire \Add0~14_combout ;
wire \counter~20_combout ;
wire \counter[7]~8_combout ;
wire \Add3~13 ;
wire \Add3~14_combout ;
wire \counter[7]~q ;
wire \Add0~15 ;
wire \Add0~16_combout ;
wire \counter[8]~7_combout ;
wire \Add3~15 ;
wire \Add3~16_combout ;
wire \counter[9]~18_combout ;
wire \counter[8]~q ;
wire \Add0~17 ;
wire \Add0~18_combout ;
wire \counter[9]~6_combout ;
wire \Add3~17 ;
wire \Add3~18_combout ;
wire \counter[9]~q ;
wire \Add0~19 ;
wire \Add0~20_combout ;
wire \counter[10]~5_combout ;
wire \Add3~19 ;
wire \Add3~20_combout ;
wire \counter[10]~q ;
wire \Add0~21 ;
wire \Add0~22_combout ;
wire \counter[11]~4_combout ;
wire \Add3~21 ;
wire \Add3~22_combout ;
wire \counter[11]~q ;
wire \Add0~23 ;
wire \Add0~24_combout ;
wire \counter[12]~3_combout ;
wire \Add3~23 ;
wire \Add3~24_combout ;
wire \counter[12]~q ;
wire \Add0~25 ;
wire \Add0~26_combout ;
wire \counter[13]~2_combout ;
wire \Add3~25 ;
wire \Add3~26_combout ;
wire \counter[13]~q ;
wire \Add0~27 ;
wire \Add0~28_combout ;
wire \counter[14]~1_combout ;
wire \Add3~27 ;
wire \Add3~28_combout ;
wire \counter[14]~q ;
wire \Add0~29 ;
wire \Add0~30_combout ;
wire \counter[15]~0_combout ;
wire \Add3~29 ;
wire \Add3~30_combout ;
wire \counter[15]~q ;
wire \Equal10~0_combout ;
wire \Equal10~1_combout ;
wire \Equal10~2_combout ;
wire \Equal10~3_combout ;
wire \Equal10~4_combout ;
wire \state~68_combout ;
wire \state~69_combout ;
wire \state.0000~q ;
wire \state~48_combout ;
wire \state~65_combout ;
wire \state~66_combout ;
wire \state.GET_EXTRA~2_combout ;
wire \state.GET_EXTRA~q ;
wire \state~73_combout ;
wire \state.GET_SIZE1~q ;
wire \state~74_combout ;
wire \state.GET_SIZE2~q ;
wire \state~75_combout ;
wire \state.GET_ADDR1~q ;
wire \state~76_combout ;
wire \state.GET_ADDR2~q ;
wire \state~77_combout ;
wire \state.GET_ADDR3~q ;
wire \state~63_combout ;
wire \state.GET_ADDR4~q ;
wire \state~72_combout ;
wire \Selector1~0_combout ;
wire \in_ready_0~4_combout ;
wire \state~81_combout ;
wire \state.GET_WRITE_DATA~q ;
wire \state~64_combout ;
wire \state~67_combout ;
wire \state.WRITE_WAIT~q ;
wire \out_data[0]~5_combout ;
wire \WideOr14~0_combout ;
wire \current_byte[1]~1_combout ;
wire \current_byte[1]~2_combout ;
wire \out_data[0]~6_combout ;
wire \current_byte[0]~3_combout ;
wire \current_byte[0]~4_combout ;
wire \current_byte[0]~q ;
wire \Selector70~0_combout ;
wire \Selector70~1_combout ;
wire \current_byte[1]~q ;
wire \Selector82~0_combout ;
wire \out_endofpacket~0_combout ;
wire \read_data_buffer[0]~q ;
wire \out_data[0]~0_combout ;
wire \out_data[0]~1_combout ;
wire \Selector80~0_combout ;
wire \Selector80~1_combout ;
wire \out_data[0]~2_combout ;
wire \out_data[0]~3_combout ;
wire \Selector80~2_combout ;
wire \WideOr14~1_combout ;
wire \out_data[0]~8_combout ;
wire \out_data[0]~9_combout ;
wire \out_data[0]~10_combout ;
wire \Selector72~0_combout ;
wire \Selector38~0_combout ;
wire \first_trans~q ;
wire \Selector72~2_combout ;
wire \Selector72~3_combout ;
wire \read_data_buffer[2]~q ;
wire \command[2]~q ;
wire \Selector78~0_combout ;
wire \Selector78~1_combout ;
wire \Selector78~2_combout ;
wire \read_data_buffer[1]~q ;
wire \Selector79~0_combout ;
wire \Selector79~1_combout ;
wire \Selector79~2_combout ;
wire \read_data_buffer[5]~q ;
wire \Selector75~0_combout ;
wire \Selector75~1_combout ;
wire \Selector75~2_combout ;
wire \read_data_buffer[7]~q ;
wire \Selector73~0_combout ;
wire \Selector73~1_combout ;
wire \Selector73~2_combout ;
wire \Selector73~3_combout ;
wire \WideOr14~2_combout ;
wire \Selector73~4_combout ;
wire \Selector73~5_combout ;
wire \read_data_buffer[6]~q ;
wire \Selector74~0_combout ;
wire \Selector74~1_combout ;
wire \Selector74~2_combout ;
wire \read_data_buffer[4]~q ;
wire \Selector76~0_combout ;
wire \Selector76~1_combout ;
wire \Selector76~2_combout ;
wire \read_data_buffer[3]~q ;
wire \Selector77~0_combout ;
wire \Selector77~1_combout ;
wire \Selector77~2_combout ;
wire \Selector0~0_combout ;
wire \Selector0~1_combout ;
wire \Selector0~2_combout ;
wire \Add2~1 ;
wire \Add2~3 ;
wire \Add2~5 ;
wire \Add2~7 ;
wire \Add2~9 ;
wire \Add2~10_combout ;
wire \Selector64~0_combout ;
wire \address[9]~3_combout ;
wire \address[9]~4_combout ;
wire \address[4]~6_combout ;
wire \Add2~8_combout ;
wire \Selector65~0_combout ;
wire \Add2~6_combout ;
wire \Selector66~0_combout ;
wire \Add2~4_combout ;
wire \Selector67~0_combout ;
wire \Add2~11 ;
wire \Add2~13 ;
wire \Add2~14_combout ;
wire \Selector62~0_combout ;
wire \address[9]~5_combout ;
wire \Add2~2_combout ;
wire \Selector68~0_combout ;
wire \Add2~12_combout ;
wire \Selector63~0_combout ;
wire \Selector81~0_combout ;
wire \in_ready_0~2_combout ;
wire \in_ready_0~3_combout ;
wire \in_ready_0~5_combout ;
wire \Selector83~0_combout ;
wire \Selector83~1_combout ;
wire \Add2~0_combout ;
wire \Selector69~0_combout ;
wire \writedata[3]~0_combout ;


dffeas out_endofpacket(
	.clk(clk),
	.d(\out_endofpacket~0_combout ),
	.asdata(\Equal10~4_combout ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.READ_SEND_ISSUE~q ),
	.ena(vcc),
	.q(out_endofpacket1),
	.prn(vcc));
defparam out_endofpacket.is_wysiwyg = "true";
defparam out_endofpacket.power_up = "low";

dffeas \out_data[0] (
	.clk(clk),
	.d(\Selector80~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_data[0]~10_combout ),
	.q(out_data_0),
	.prn(vcc));
defparam \out_data[0] .is_wysiwyg = "true";
defparam \out_data[0] .power_up = "low";

dffeas out_startofpacket(
	.clk(clk),
	.d(\Selector72~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_startofpacket1),
	.prn(vcc));
defparam out_startofpacket.is_wysiwyg = "true";
defparam out_startofpacket.power_up = "low";

dffeas \out_data[2] (
	.clk(clk),
	.d(\Selector78~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_data[0]~10_combout ),
	.q(out_data_2),
	.prn(vcc));
defparam \out_data[2] .is_wysiwyg = "true";
defparam \out_data[2] .power_up = "low";

dffeas \out_data[1] (
	.clk(clk),
	.d(\Selector79~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_data[0]~10_combout ),
	.q(out_data_1),
	.prn(vcc));
defparam \out_data[1] .is_wysiwyg = "true";
defparam \out_data[1] .power_up = "low";

dffeas \out_data[5] (
	.clk(clk),
	.d(\Selector75~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_data[0]~10_combout ),
	.q(out_data_5),
	.prn(vcc));
defparam \out_data[5] .is_wysiwyg = "true";
defparam \out_data[5] .power_up = "low";

dffeas \out_data[7] (
	.clk(clk),
	.d(\Selector73~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_data_7),
	.prn(vcc));
defparam \out_data[7] .is_wysiwyg = "true";
defparam \out_data[7] .power_up = "low";

dffeas \out_data[6] (
	.clk(clk),
	.d(\Selector74~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_data[0]~10_combout ),
	.q(out_data_6),
	.prn(vcc));
defparam \out_data[6] .is_wysiwyg = "true";
defparam \out_data[6] .power_up = "low";

dffeas \out_data[4] (
	.clk(clk),
	.d(\Selector76~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_data[0]~10_combout ),
	.q(out_data_4),
	.prn(vcc));
defparam \out_data[4] .is_wysiwyg = "true";
defparam \out_data[4] .power_up = "low";

dffeas \out_data[3] (
	.clk(clk),
	.d(\Selector77~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_data[0]~10_combout ),
	.q(out_data_3),
	.prn(vcc));
defparam \out_data[3] .is_wysiwyg = "true";
defparam \out_data[3] .power_up = "low";

dffeas out_valid(
	.clk(clk),
	.d(\Selector0~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_valid1),
	.prn(vcc));
defparam out_valid.is_wysiwyg = "true";
defparam out_valid.power_up = "low";

dffeas \address[7] (
	.clk(clk),
	.d(\Selector64~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address[4]~6_combout ),
	.q(address_7),
	.prn(vcc));
defparam \address[7] .is_wysiwyg = "true";
defparam \address[7] .power_up = "low";

dffeas \address[6] (
	.clk(clk),
	.d(\Selector65~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address[4]~6_combout ),
	.q(address_6),
	.prn(vcc));
defparam \address[6] .is_wysiwyg = "true";
defparam \address[6] .power_up = "low";

dffeas \address[5] (
	.clk(clk),
	.d(\Selector66~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address[4]~6_combout ),
	.q(address_5),
	.prn(vcc));
defparam \address[5] .is_wysiwyg = "true";
defparam \address[5] .power_up = "low";

dffeas \address[4] (
	.clk(clk),
	.d(\Selector67~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address[4]~6_combout ),
	.q(address_4),
	.prn(vcc));
defparam \address[4] .is_wysiwyg = "true";
defparam \address[4] .power_up = "low";

dffeas \address[9] (
	.clk(clk),
	.d(\Selector62~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address[9]~5_combout ),
	.q(address_9),
	.prn(vcc));
defparam \address[9] .is_wysiwyg = "true";
defparam \address[9] .power_up = "low";

dffeas \address[3] (
	.clk(clk),
	.d(\Selector68~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address[4]~6_combout ),
	.q(address_3),
	.prn(vcc));
defparam \address[3] .is_wysiwyg = "true";
defparam \address[3] .power_up = "low";

dffeas \address[8] (
	.clk(clk),
	.d(\Selector63~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address[9]~5_combout ),
	.q(address_8),
	.prn(vcc));
defparam \address[8] .is_wysiwyg = "true";
defparam \address[8] .power_up = "low";

dffeas write(
	.clk(clk),
	.d(\Selector81~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(write1),
	.prn(vcc));
defparam write.is_wysiwyg = "true";
defparam write.power_up = "low";

dffeas in_ready_0(
	.clk(clk),
	.d(\in_ready_0~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(in_ready_01),
	.prn(vcc));
defparam in_ready_0.is_wysiwyg = "true";
defparam in_ready_0.power_up = "low";

fiftyfivenm_lcell_comb \enable~0 (
	.dataa(out_valid3),
	.datab(in_ready_01),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(enable1),
	.cout());
defparam \enable~0 .lut_mask = 16'hEEEE;
defparam \enable~0 .sum_lutc_input = "datac";

dffeas read(
	.clk(clk),
	.d(\Selector83~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read1),
	.prn(vcc));
defparam read.is_wysiwyg = "true";
defparam read.power_up = "low";

dffeas \address[2] (
	.clk(clk),
	.d(\Selector69~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\address[4]~6_combout ),
	.q(address_2),
	.prn(vcc));
defparam \address[2] .is_wysiwyg = "true";
defparam \address[2] .power_up = "low";

dffeas \writedata[0] (
	.clk(clk),
	.d(in_data[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\writedata[3]~0_combout ),
	.q(writedata_0),
	.prn(vcc));
defparam \writedata[0] .is_wysiwyg = "true";
defparam \writedata[0] .power_up = "low";

dffeas \writedata[2] (
	.clk(clk),
	.d(in_data[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\writedata[3]~0_combout ),
	.q(writedata_2),
	.prn(vcc));
defparam \writedata[2] .is_wysiwyg = "true";
defparam \writedata[2] .power_up = "low";

dffeas \writedata[1] (
	.clk(clk),
	.d(in_data[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\writedata[3]~0_combout ),
	.q(writedata_1),
	.prn(vcc));
defparam \writedata[1] .is_wysiwyg = "true";
defparam \writedata[1] .power_up = "low";

dffeas \writedata[3] (
	.clk(clk),
	.d(in_data[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\writedata[3]~0_combout ),
	.q(writedata_3),
	.prn(vcc));
defparam \writedata[3] .is_wysiwyg = "true";
defparam \writedata[3] .power_up = "low";

fiftyfivenm_lcell_comb \enable~1 (
	.dataa(out_channel_0),
	.datab(out_channel_7),
	.datac(out_channel_6),
	.datad(out_channel_5),
	.cin(gnd),
	.combout(\enable~1_combout ),
	.cout());
defparam \enable~1 .lut_mask = 16'h7FFF;
defparam \enable~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \enable~2 (
	.dataa(out_channel_4),
	.datab(out_channel_3),
	.datac(out_channel_2),
	.datad(out_channel_1),
	.cin(gnd),
	.combout(\enable~2_combout ),
	.cout());
defparam \enable~2 .lut_mask = 16'h7FFF;
defparam \enable~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \enable~3 (
	.dataa(\enable~1_combout ),
	.datab(\enable~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\enable~3_combout ),
	.cout());
defparam \enable~3 .lut_mask = 16'hEEEE;
defparam \enable~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb enable(
	.dataa(out_valid2),
	.datab(enable1),
	.datac(\enable~3_combout ),
	.datad(received_channel),
	.cin(gnd),
	.combout(\enable~combout ),
	.cout());
defparam enable.lut_mask = 16'hFEFF;
defparam enable.sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \always1~0 (
	.dataa(\enable~combout ),
	.datab(out_startofpacket2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\always1~0_combout ),
	.cout());
defparam \always1~0 .lut_mask = 16'hEEEE;
defparam \always1~0 .sum_lutc_input = "datac";

dffeas \command[7] (
	.clk(clk),
	.d(in_data[7]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(\command[7]~q ),
	.prn(vcc));
defparam \command[7] .is_wysiwyg = "true";
defparam \command[7] .power_up = "low";

dffeas \command[6] (
	.clk(clk),
	.d(in_data[6]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(\command[6]~q ),
	.prn(vcc));
defparam \command[6] .is_wysiwyg = "true";
defparam \command[6] .power_up = "low";

dffeas \command[5] (
	.clk(clk),
	.d(in_data[5]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(\command[5]~q ),
	.prn(vcc));
defparam \command[5] .is_wysiwyg = "true";
defparam \command[5] .power_up = "low";

dffeas \command[3] (
	.clk(clk),
	.d(in_data[3]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(\command[3]~q ),
	.prn(vcc));
defparam \command[3] .is_wysiwyg = "true";
defparam \command[3] .power_up = "low";

fiftyfivenm_lcell_comb \Equal2~0 (
	.dataa(\command[7]~q ),
	.datab(\command[6]~q ),
	.datac(\command[5]~q ),
	.datad(\command[3]~q ),
	.cin(gnd),
	.combout(\Equal2~0_combout ),
	.cout());
defparam \Equal2~0 .lut_mask = 16'h7FFF;
defparam \Equal2~0 .sum_lutc_input = "datac";

dffeas \command[0] (
	.clk(clk),
	.d(in_data[0]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(\command[0]~q ),
	.prn(vcc));
defparam \command[0] .is_wysiwyg = "true";
defparam \command[0] .power_up = "low";

dffeas \command[1] (
	.clk(clk),
	.d(in_data[1]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(\command[1]~q ),
	.prn(vcc));
defparam \command[1] .is_wysiwyg = "true";
defparam \command[1] .power_up = "low";

fiftyfivenm_lcell_comb \Equal2~1 (
	.dataa(\Equal2~0_combout ),
	.datab(gnd),
	.datac(\command[0]~q ),
	.datad(\command[1]~q ),
	.cin(gnd),
	.combout(\Equal2~1_combout ),
	.cout());
defparam \Equal2~1 .lut_mask = 16'hAFFF;
defparam \Equal2~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector72~1 (
	.dataa(\state.GET_ADDR4~q ),
	.datab(\enable~combout ),
	.datac(gnd),
	.datad(\Equal2~1_combout ),
	.cin(gnd),
	.combout(\Selector72~1_combout ),
	.cout());
defparam \Selector72~1 .lut_mask = 16'hEEFF;
defparam \Selector72~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector39~0 (
	.dataa(\state.GET_WRITE_DATA~q ),
	.datab(\last_trans~q ),
	.datac(out_endofpacket2),
	.datad(\state.GET_ADDR1~q ),
	.cin(gnd),
	.combout(\Selector39~0_combout ),
	.cout());
defparam \Selector39~0 .lut_mask = 16'hFEFF;
defparam \Selector39~0 .sum_lutc_input = "datac";

dffeas last_trans(
	.clk(clk),
	.d(\Selector39~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\last_trans~q ),
	.prn(vcc));
defparam last_trans.is_wysiwyg = "true";
defparam last_trans.power_up = "low";

fiftyfivenm_lcell_comb \state~59 (
	.dataa(\Selector72~1_combout ),
	.datab(\state.WRITE_WAIT~q ),
	.datac(\last_trans~q ),
	.datad(av_waitrequest),
	.cin(gnd),
	.combout(\state~59_combout ),
	.cout());
defparam \state~59 .lut_mask = 16'hFEFF;
defparam \state~59 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \state~79 (
	.dataa(\current_byte[1]~q ),
	.datab(\current_byte[0]~q ),
	.datac(in_ready),
	.datad(gnd),
	.cin(gnd),
	.combout(\state~79_combout ),
	.cout());
defparam \state~79 .lut_mask = 16'hFEFE;
defparam \state~79 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \state~60 (
	.dataa(\state~59_combout ),
	.datab(\state.RETURN_PACKET~q ),
	.datac(\state~79_combout ),
	.datad(\always1~0_combout ),
	.cin(gnd),
	.combout(\state~60_combout ),
	.cout());
defparam \state~60 .lut_mask = 16'hEFFF;
defparam \state~60 .sum_lutc_input = "datac";

dffeas \state.RETURN_PACKET (
	.clk(clk),
	.d(\state~60_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.RETURN_PACKET~q ),
	.prn(vcc));
defparam \state.RETURN_PACKET .is_wysiwyg = "true";
defparam \state.RETURN_PACKET .power_up = "low";

fiftyfivenm_lcell_comb \Add0~0 (
	.dataa(\counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout(\Add0~1 ));
defparam \Add0~0 .lut_mask = 16'h55AA;
defparam \Add0~0 .sum_lutc_input = "datac";

dffeas \command[4] (
	.clk(clk),
	.d(in_data[4]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(\command[4]~q ),
	.prn(vcc));
defparam \command[4] .is_wysiwyg = "true";
defparam \command[4] .power_up = "low";

fiftyfivenm_lcell_comb \counter~16 (
	.dataa(\command[4]~q ),
	.datab(in_data[0]),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\counter~16_combout ),
	.cout());
defparam \counter~16 .lut_mask = 16'hEEEE;
defparam \counter~16 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \counter[0]~15 (
	.dataa(\Add0~0_combout ),
	.datab(\counter~16_combout ),
	.datac(gnd),
	.datad(\state.GET_WRITE_DATA~q ),
	.cin(gnd),
	.combout(\counter[0]~15_combout ),
	.cout());
defparam \counter[0]~15 .lut_mask = 16'hAACC;
defparam \counter[0]~15 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add3~0 (
	.dataa(\counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add3~0_combout ),
	.cout(\Add3~1 ));
defparam \Add3~0 .lut_mask = 16'h55AA;
defparam \Add3~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data[0]~7 (
	.dataa(\current_byte[1]~q ),
	.datab(\current_byte[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_data[0]~7_combout ),
	.cout());
defparam \out_data[0]~7 .lut_mask = 16'hEEEE;
defparam \out_data[0]~7 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \state~61 (
	.dataa(in_ready),
	.datab(\state.READ_SEND_WAIT~q ),
	.datac(\out_data[0]~7_combout ),
	.datad(\Equal10~4_combout ),
	.cin(gnd),
	.combout(\state~61_combout ),
	.cout());
defparam \state~61 .lut_mask = 16'hEFFF;
defparam \state~61 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \address[9]~2 (
	.dataa(in_ready),
	.datab(\out_data[0]~7_combout ),
	.datac(\state.READ_SEND_WAIT~q ),
	.datad(\Equal10~4_combout ),
	.cin(gnd),
	.combout(\address[9]~2_combout ),
	.cout());
defparam \address[9]~2 .lut_mask = 16'hFEFF;
defparam \address[9]~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \state~71 (
	.dataa(\state.GET_ADDR4~q ),
	.datab(\command[4]~q ),
	.datac(\Equal2~1_combout ),
	.datad(\enable~combout ),
	.cin(gnd),
	.combout(\state~71_combout ),
	.cout());
defparam \state~71 .lut_mask = 16'hFFFE;
defparam \state~71 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \state~80 (
	.dataa(\enable~combout ),
	.datab(out_startofpacket2),
	.datac(\address[9]~2_combout ),
	.datad(\state~71_combout ),
	.cin(gnd),
	.combout(\state~80_combout ),
	.cout());
defparam \state~80 .lut_mask = 16'hFFF7;
defparam \state~80 .sum_lutc_input = "datac";

dffeas \state.READ_ASSERT (
	.clk(clk),
	.d(\state~80_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.READ_ASSERT~q ),
	.prn(vcc));
defparam \state.READ_ASSERT .is_wysiwyg = "true";
defparam \state.READ_ASSERT .power_up = "low";

fiftyfivenm_lcell_comb \state~49 (
	.dataa(\state.RETURN_PACKET~q ),
	.datab(\state.WRITE_WAIT~q ),
	.datac(\state.READ_SEND_WAIT~q ),
	.datad(\out_data~4_combout ),
	.cin(gnd),
	.combout(\state~49_combout ),
	.cout());
defparam \state~49 .lut_mask = 16'hFFFE;
defparam \state~49 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \state~58 (
	.dataa(\state.READ_DATA_WAIT~q ),
	.datab(\state.READ_CMD_WAIT~q ),
	.datac(av_waitrequest),
	.datad(WideOr1),
	.cin(gnd),
	.combout(\state~58_combout ),
	.cout());
defparam \state~58 .lut_mask = 16'hEFFF;
defparam \state~58 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \state~78 (
	.dataa(\enable~combout ),
	.datab(out_startofpacket2),
	.datac(\state~58_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\state~78_combout ),
	.cout());
defparam \state~78 .lut_mask = 16'hF7F7;
defparam \state~78 .sum_lutc_input = "datac";

dffeas \state.READ_DATA_WAIT (
	.clk(clk),
	.d(\state~78_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.READ_DATA_WAIT~q ),
	.prn(vcc));
defparam \state.READ_DATA_WAIT .is_wysiwyg = "true";
defparam \state.READ_DATA_WAIT .power_up = "low";

fiftyfivenm_lcell_comb \current_byte[1]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\state.RETURN_PACKET~q ),
	.datad(\state.READ_SEND_WAIT~q ),
	.cin(gnd),
	.combout(\current_byte[1]~0_combout ),
	.cout());
defparam \current_byte[1]~0 .lut_mask = 16'h0FFF;
defparam \current_byte[1]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \state~50 (
	.dataa(WideOr1),
	.datab(\state.READ_DATA_WAIT~q ),
	.datac(in_ready),
	.datad(\current_byte[1]~0_combout ),
	.cin(gnd),
	.combout(\state~50_combout ),
	.cout());
defparam \state~50 .lut_mask = 16'hB8FF;
defparam \state~50 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \state~51 (
	.dataa(\state.READ_CMD_WAIT~q ),
	.datab(\state.WRITE_WAIT~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\state~51_combout ),
	.cout());
defparam \state~51 .lut_mask = 16'hEEEE;
defparam \state~51 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \state~52 (
	.dataa(\state~49_combout ),
	.datab(\state~50_combout ),
	.datac(\state~51_combout ),
	.datad(av_waitrequest),
	.cin(gnd),
	.combout(\state~52_combout ),
	.cout());
defparam \state~52 .lut_mask = 16'hFEFF;
defparam \state~52 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \state~53 (
	.dataa(\state.READ_CMD_WAIT~q ),
	.datab(WideOr1),
	.datac(\state.READ_SEND_ISSUE~q ),
	.datad(\state.READ_ASSERT~q ),
	.cin(gnd),
	.combout(\state~53_combout ),
	.cout());
defparam \state~53 .lut_mask = 16'h7FFF;
defparam \state~53 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \write~0 (
	.dataa(out_endofpacket2),
	.datab(\current_byte[1]~q ),
	.datac(\current_byte[0]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\write~0_combout ),
	.cout());
defparam \write~0 .lut_mask = 16'hFEFE;
defparam \write~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \in_ready_0~0 (
	.dataa(\state.GET_EXTRA~q ),
	.datab(\state.GET_SIZE1~q ),
	.datac(\state.GET_SIZE2~q ),
	.datad(\state.GET_ADDR1~q ),
	.cin(gnd),
	.combout(\in_ready_0~0_combout ),
	.cout());
defparam \in_ready_0~0 .lut_mask = 16'h7FFF;
defparam \in_ready_0~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \in_ready_0~1 (
	.dataa(\in_ready_0~0_combout ),
	.datab(gnd),
	.datac(\state.GET_ADDR2~q ),
	.datad(\state.GET_ADDR3~q ),
	.cin(gnd),
	.combout(\in_ready_0~1_combout ),
	.cout());
defparam \in_ready_0~1 .lut_mask = 16'hAFFF;
defparam \in_ready_0~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \state~54 (
	.dataa(\state.GET_WRITE_DATA~q ),
	.datab(\write~0_combout ),
	.datac(\state.GET_ADDR4~q ),
	.datad(\in_ready_0~1_combout ),
	.cin(gnd),
	.combout(\state~54_combout ),
	.cout());
defparam \state~54 .lut_mask = 16'hFF7F;
defparam \state~54 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \state~55 (
	.dataa(\enable~combout ),
	.datab(\state.0000~q ),
	.datac(out_startofpacket2),
	.datad(\state~54_combout ),
	.cin(gnd),
	.combout(\state~55_combout ),
	.cout());
defparam \state~55 .lut_mask = 16'hFEFF;
defparam \state~55 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \state~56 (
	.dataa(\state~48_combout ),
	.datab(\state~52_combout ),
	.datac(\state~53_combout ),
	.datad(\state~55_combout ),
	.cin(gnd),
	.combout(\state~56_combout ),
	.cout());
defparam \state~56 .lut_mask = 16'hFFEF;
defparam \state~56 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \state~57 (
	.dataa(\state.READ_CMD_WAIT~q ),
	.datab(\state.READ_ASSERT~q ),
	.datac(\state~56_combout ),
	.datad(\always1~0_combout ),
	.cin(gnd),
	.combout(\state~57_combout ),
	.cout());
defparam \state~57 .lut_mask = 16'hEFFF;
defparam \state~57 .sum_lutc_input = "datac";

dffeas \state.READ_CMD_WAIT (
	.clk(clk),
	.d(\state~57_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.READ_CMD_WAIT~q ),
	.prn(vcc));
defparam \state.READ_CMD_WAIT .is_wysiwyg = "true";
defparam \state.READ_CMD_WAIT .power_up = "low";

fiftyfivenm_lcell_comb \out_data~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\state.READ_CMD_WAIT~q ),
	.datad(\state.READ_DATA_WAIT~q ),
	.cin(gnd),
	.combout(\out_data~4_combout ),
	.cout());
defparam \out_data~4 .lut_mask = 16'hFFF0;
defparam \out_data~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \state~62 (
	.dataa(\state~61_combout ),
	.datab(WideOr1),
	.datac(\out_data~4_combout ),
	.datad(\always1~0_combout ),
	.cin(gnd),
	.combout(\state~62_combout ),
	.cout());
defparam \state~62 .lut_mask = 16'hFEFF;
defparam \state~62 .sum_lutc_input = "datac";

dffeas \state.READ_SEND_ISSUE (
	.clk(clk),
	.d(\state~62_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.READ_SEND_ISSUE~q ),
	.prn(vcc));
defparam \state.READ_SEND_ISSUE .is_wysiwyg = "true";
defparam \state.READ_SEND_ISSUE .power_up = "low";

fiftyfivenm_lcell_comb \state~70 (
	.dataa(\state.READ_SEND_ISSUE~q ),
	.datab(\state.READ_SEND_WAIT~q ),
	.datac(\always1~0_combout ),
	.datad(\state~56_combout ),
	.cin(gnd),
	.combout(\state~70_combout ),
	.cout());
defparam \state~70 .lut_mask = 16'hEFFF;
defparam \state~70 .sum_lutc_input = "datac";

dffeas \state.READ_SEND_WAIT (
	.clk(clk),
	.d(\state~70_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.READ_SEND_WAIT~q ),
	.prn(vcc));
defparam \state.READ_SEND_WAIT .is_wysiwyg = "true";
defparam \state.READ_SEND_WAIT .power_up = "low";

fiftyfivenm_lcell_comb \counter[9]~17 (
	.dataa(in_ready),
	.datab(\enable~combout ),
	.datac(\state.GET_WRITE_DATA~q ),
	.datad(\state.READ_SEND_WAIT~q ),
	.cin(gnd),
	.combout(\counter[9]~17_combout ),
	.cout());
defparam \counter[9]~17 .lut_mask = 16'hEFFF;
defparam \counter[9]~17 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \counter[4]~19 (
	.dataa(\state.READ_SEND_WAIT~q ),
	.datab(\state.GET_WRITE_DATA~q ),
	.datac(\state.GET_SIZE2~q ),
	.datad(\counter[9]~17_combout ),
	.cin(gnd),
	.combout(\counter[4]~19_combout ),
	.cout());
defparam \counter[4]~19 .lut_mask = 16'hFFFE;
defparam \counter[4]~19 .sum_lutc_input = "datac";

dffeas \counter[0] (
	.clk(clk),
	.d(\counter[0]~15_combout ),
	.asdata(\Add3~0_combout ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.READ_SEND_WAIT~q ),
	.ena(\counter[4]~19_combout ),
	.q(\counter[0]~q ),
	.prn(vcc));
defparam \counter[0] .is_wysiwyg = "true";
defparam \counter[0] .power_up = "low";

fiftyfivenm_lcell_comb \Add0~2 (
	.dataa(\counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~1 ),
	.combout(\Add0~2_combout ),
	.cout(\Add0~3 ));
defparam \Add0~2 .lut_mask = 16'h5A5F;
defparam \Add0~2 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \counter~26 (
	.dataa(\command[4]~q ),
	.datab(in_data[1]),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\counter~26_combout ),
	.cout());
defparam \counter~26 .lut_mask = 16'hEEEE;
defparam \counter~26 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \counter[1]~14 (
	.dataa(\Add0~2_combout ),
	.datab(\counter~26_combout ),
	.datac(gnd),
	.datad(\state.GET_WRITE_DATA~q ),
	.cin(gnd),
	.combout(\counter[1]~14_combout ),
	.cout());
defparam \counter[1]~14 .lut_mask = 16'hAACC;
defparam \counter[1]~14 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add3~2 (
	.dataa(\counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~1 ),
	.combout(\Add3~2_combout ),
	.cout(\Add3~3 ));
defparam \Add3~2 .lut_mask = 16'h5A5F;
defparam \Add3~2 .sum_lutc_input = "cin";

dffeas \counter[1] (
	.clk(clk),
	.d(\counter[1]~14_combout ),
	.asdata(\Add3~2_combout ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.READ_SEND_WAIT~q ),
	.ena(\counter[4]~19_combout ),
	.q(\counter[1]~q ),
	.prn(vcc));
defparam \counter[1] .is_wysiwyg = "true";
defparam \counter[1] .power_up = "low";

fiftyfivenm_lcell_comb \Add0~4 (
	.dataa(\counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~3 ),
	.combout(\Add0~4_combout ),
	.cout(\Add0~5 ));
defparam \Add0~4 .lut_mask = 16'h5AAF;
defparam \Add0~4 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \counter~25 (
	.dataa(\command[4]~q ),
	.datab(in_data[2]),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\counter~25_combout ),
	.cout());
defparam \counter~25 .lut_mask = 16'hEEEE;
defparam \counter~25 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \counter[2]~13 (
	.dataa(\Add0~4_combout ),
	.datab(\counter~25_combout ),
	.datac(gnd),
	.datad(\state.GET_WRITE_DATA~q ),
	.cin(gnd),
	.combout(\counter[2]~13_combout ),
	.cout());
defparam \counter[2]~13 .lut_mask = 16'hAACC;
defparam \counter[2]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add3~4 (
	.dataa(\counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~3 ),
	.combout(\Add3~4_combout ),
	.cout(\Add3~5 ));
defparam \Add3~4 .lut_mask = 16'h5AAF;
defparam \Add3~4 .sum_lutc_input = "cin";

dffeas \counter[2] (
	.clk(clk),
	.d(\counter[2]~13_combout ),
	.asdata(\Add3~4_combout ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.READ_SEND_WAIT~q ),
	.ena(\counter[4]~19_combout ),
	.q(\counter[2]~q ),
	.prn(vcc));
defparam \counter[2] .is_wysiwyg = "true";
defparam \counter[2] .power_up = "low";

fiftyfivenm_lcell_comb \Add0~6 (
	.dataa(\counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~5 ),
	.combout(\Add0~6_combout ),
	.cout(\Add0~7 ));
defparam \Add0~6 .lut_mask = 16'h5A5F;
defparam \Add0~6 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \counter~24 (
	.dataa(\command[4]~q ),
	.datab(in_data[3]),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\counter~24_combout ),
	.cout());
defparam \counter~24 .lut_mask = 16'hEEEE;
defparam \counter~24 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \counter[3]~12 (
	.dataa(\Add0~6_combout ),
	.datab(\counter~24_combout ),
	.datac(gnd),
	.datad(\state.GET_WRITE_DATA~q ),
	.cin(gnd),
	.combout(\counter[3]~12_combout ),
	.cout());
defparam \counter[3]~12 .lut_mask = 16'hAACC;
defparam \counter[3]~12 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add3~6 (
	.dataa(\counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~5 ),
	.combout(\Add3~6_combout ),
	.cout(\Add3~7 ));
defparam \Add3~6 .lut_mask = 16'h5A5F;
defparam \Add3~6 .sum_lutc_input = "cin";

dffeas \counter[3] (
	.clk(clk),
	.d(\counter[3]~12_combout ),
	.asdata(\Add3~6_combout ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.READ_SEND_WAIT~q ),
	.ena(\counter[4]~19_combout ),
	.q(\counter[3]~q ),
	.prn(vcc));
defparam \counter[3] .is_wysiwyg = "true";
defparam \counter[3] .power_up = "low";

fiftyfivenm_lcell_comb \Add0~8 (
	.dataa(\counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~7 ),
	.combout(\Add0~8_combout ),
	.cout(\Add0~9 ));
defparam \Add0~8 .lut_mask = 16'h5AAF;
defparam \Add0~8 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \counter~23 (
	.dataa(\command[4]~q ),
	.datab(in_data[4]),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\counter~23_combout ),
	.cout());
defparam \counter~23 .lut_mask = 16'hEEEE;
defparam \counter~23 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \counter[4]~11 (
	.dataa(\Add0~8_combout ),
	.datab(\counter~23_combout ),
	.datac(gnd),
	.datad(\state.GET_WRITE_DATA~q ),
	.cin(gnd),
	.combout(\counter[4]~11_combout ),
	.cout());
defparam \counter[4]~11 .lut_mask = 16'hAACC;
defparam \counter[4]~11 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add3~8 (
	.dataa(\counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~7 ),
	.combout(\Add3~8_combout ),
	.cout(\Add3~9 ));
defparam \Add3~8 .lut_mask = 16'h5AAF;
defparam \Add3~8 .sum_lutc_input = "cin";

dffeas \counter[4] (
	.clk(clk),
	.d(\counter[4]~11_combout ),
	.asdata(\Add3~8_combout ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.READ_SEND_WAIT~q ),
	.ena(\counter[4]~19_combout ),
	.q(\counter[4]~q ),
	.prn(vcc));
defparam \counter[4] .is_wysiwyg = "true";
defparam \counter[4] .power_up = "low";

fiftyfivenm_lcell_comb \Add0~10 (
	.dataa(\counter[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~9 ),
	.combout(\Add0~10_combout ),
	.cout(\Add0~11 ));
defparam \Add0~10 .lut_mask = 16'h5A5F;
defparam \Add0~10 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \counter~22 (
	.dataa(\command[4]~q ),
	.datab(gnd),
	.datac(received_esc),
	.datad(out_payload_5),
	.cin(gnd),
	.combout(\counter~22_combout ),
	.cout());
defparam \counter~22 .lut_mask = 16'hAFFA;
defparam \counter~22 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \counter[5]~10 (
	.dataa(\Add0~10_combout ),
	.datab(\counter~22_combout ),
	.datac(gnd),
	.datad(\state.GET_WRITE_DATA~q ),
	.cin(gnd),
	.combout(\counter[5]~10_combout ),
	.cout());
defparam \counter[5]~10 .lut_mask = 16'hAACC;
defparam \counter[5]~10 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add3~10 (
	.dataa(\counter[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~9 ),
	.combout(\Add3~10_combout ),
	.cout(\Add3~11 ));
defparam \Add3~10 .lut_mask = 16'h5A5F;
defparam \Add3~10 .sum_lutc_input = "cin";

dffeas \counter[5] (
	.clk(clk),
	.d(\counter[5]~10_combout ),
	.asdata(\Add3~10_combout ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.READ_SEND_WAIT~q ),
	.ena(\counter[4]~19_combout ),
	.q(\counter[5]~q ),
	.prn(vcc));
defparam \counter[5] .is_wysiwyg = "true";
defparam \counter[5] .power_up = "low";

fiftyfivenm_lcell_comb \Add0~12 (
	.dataa(\counter[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~11 ),
	.combout(\Add0~12_combout ),
	.cout(\Add0~13 ));
defparam \Add0~12 .lut_mask = 16'h5AAF;
defparam \Add0~12 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \counter~21 (
	.dataa(\command[4]~q ),
	.datab(in_data[6]),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\counter~21_combout ),
	.cout());
defparam \counter~21 .lut_mask = 16'hEEEE;
defparam \counter~21 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \counter[6]~9 (
	.dataa(\Add0~12_combout ),
	.datab(\counter~21_combout ),
	.datac(gnd),
	.datad(\state.GET_WRITE_DATA~q ),
	.cin(gnd),
	.combout(\counter[6]~9_combout ),
	.cout());
defparam \counter[6]~9 .lut_mask = 16'hAACC;
defparam \counter[6]~9 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add3~12 (
	.dataa(\counter[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~11 ),
	.combout(\Add3~12_combout ),
	.cout(\Add3~13 ));
defparam \Add3~12 .lut_mask = 16'h5AAF;
defparam \Add3~12 .sum_lutc_input = "cin";

dffeas \counter[6] (
	.clk(clk),
	.d(\counter[6]~9_combout ),
	.asdata(\Add3~12_combout ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.READ_SEND_WAIT~q ),
	.ena(\counter[4]~19_combout ),
	.q(\counter[6]~q ),
	.prn(vcc));
defparam \counter[6] .is_wysiwyg = "true";
defparam \counter[6] .power_up = "low";

fiftyfivenm_lcell_comb \Add0~14 (
	.dataa(\counter[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~13 ),
	.combout(\Add0~14_combout ),
	.cout(\Add0~15 ));
defparam \Add0~14 .lut_mask = 16'h5A5F;
defparam \Add0~14 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \counter~20 (
	.dataa(\command[4]~q ),
	.datab(in_data[7]),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\counter~20_combout ),
	.cout());
defparam \counter~20 .lut_mask = 16'hEEEE;
defparam \counter~20 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \counter[7]~8 (
	.dataa(\Add0~14_combout ),
	.datab(\counter~20_combout ),
	.datac(gnd),
	.datad(\state.GET_WRITE_DATA~q ),
	.cin(gnd),
	.combout(\counter[7]~8_combout ),
	.cout());
defparam \counter[7]~8 .lut_mask = 16'hAACC;
defparam \counter[7]~8 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add3~14 (
	.dataa(\counter[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~13 ),
	.combout(\Add3~14_combout ),
	.cout(\Add3~15 ));
defparam \Add3~14 .lut_mask = 16'h5A5F;
defparam \Add3~14 .sum_lutc_input = "cin";

dffeas \counter[7] (
	.clk(clk),
	.d(\counter[7]~8_combout ),
	.asdata(\Add3~14_combout ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.READ_SEND_WAIT~q ),
	.ena(\counter[4]~19_combout ),
	.q(\counter[7]~q ),
	.prn(vcc));
defparam \counter[7] .is_wysiwyg = "true";
defparam \counter[7] .power_up = "low";

fiftyfivenm_lcell_comb \Add0~16 (
	.dataa(\counter[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~15 ),
	.combout(\Add0~16_combout ),
	.cout(\Add0~17 ));
defparam \Add0~16 .lut_mask = 16'h5AAF;
defparam \Add0~16 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \counter[8]~7 (
	.dataa(\Add0~16_combout ),
	.datab(\counter~16_combout ),
	.datac(gnd),
	.datad(\state.GET_WRITE_DATA~q ),
	.cin(gnd),
	.combout(\counter[8]~7_combout ),
	.cout());
defparam \counter[8]~7 .lut_mask = 16'hAACC;
defparam \counter[8]~7 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add3~16 (
	.dataa(\counter[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~15 ),
	.combout(\Add3~16_combout ),
	.cout(\Add3~17 ));
defparam \Add3~16 .lut_mask = 16'h5AAF;
defparam \Add3~16 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \counter[9]~18 (
	.dataa(\state.READ_SEND_WAIT~q ),
	.datab(\state.GET_WRITE_DATA~q ),
	.datac(\state.GET_SIZE1~q ),
	.datad(\counter[9]~17_combout ),
	.cin(gnd),
	.combout(\counter[9]~18_combout ),
	.cout());
defparam \counter[9]~18 .lut_mask = 16'hFFFE;
defparam \counter[9]~18 .sum_lutc_input = "datac";

dffeas \counter[8] (
	.clk(clk),
	.d(\counter[8]~7_combout ),
	.asdata(\Add3~16_combout ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.READ_SEND_WAIT~q ),
	.ena(\counter[9]~18_combout ),
	.q(\counter[8]~q ),
	.prn(vcc));
defparam \counter[8] .is_wysiwyg = "true";
defparam \counter[8] .power_up = "low";

fiftyfivenm_lcell_comb \Add0~18 (
	.dataa(\counter[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~17 ),
	.combout(\Add0~18_combout ),
	.cout(\Add0~19 ));
defparam \Add0~18 .lut_mask = 16'h5A5F;
defparam \Add0~18 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \counter[9]~6 (
	.dataa(\Add0~18_combout ),
	.datab(\counter~26_combout ),
	.datac(gnd),
	.datad(\state.GET_WRITE_DATA~q ),
	.cin(gnd),
	.combout(\counter[9]~6_combout ),
	.cout());
defparam \counter[9]~6 .lut_mask = 16'hAACC;
defparam \counter[9]~6 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add3~18 (
	.dataa(\counter[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~17 ),
	.combout(\Add3~18_combout ),
	.cout(\Add3~19 ));
defparam \Add3~18 .lut_mask = 16'h5A5F;
defparam \Add3~18 .sum_lutc_input = "cin";

dffeas \counter[9] (
	.clk(clk),
	.d(\counter[9]~6_combout ),
	.asdata(\Add3~18_combout ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.READ_SEND_WAIT~q ),
	.ena(\counter[9]~18_combout ),
	.q(\counter[9]~q ),
	.prn(vcc));
defparam \counter[9] .is_wysiwyg = "true";
defparam \counter[9] .power_up = "low";

fiftyfivenm_lcell_comb \Add0~20 (
	.dataa(\counter[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~19 ),
	.combout(\Add0~20_combout ),
	.cout(\Add0~21 ));
defparam \Add0~20 .lut_mask = 16'h5AAF;
defparam \Add0~20 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \counter[10]~5 (
	.dataa(\Add0~20_combout ),
	.datab(\counter~25_combout ),
	.datac(gnd),
	.datad(\state.GET_WRITE_DATA~q ),
	.cin(gnd),
	.combout(\counter[10]~5_combout ),
	.cout());
defparam \counter[10]~5 .lut_mask = 16'hAACC;
defparam \counter[10]~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add3~20 (
	.dataa(\counter[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~19 ),
	.combout(\Add3~20_combout ),
	.cout(\Add3~21 ));
defparam \Add3~20 .lut_mask = 16'h5AAF;
defparam \Add3~20 .sum_lutc_input = "cin";

dffeas \counter[10] (
	.clk(clk),
	.d(\counter[10]~5_combout ),
	.asdata(\Add3~20_combout ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.READ_SEND_WAIT~q ),
	.ena(\counter[9]~18_combout ),
	.q(\counter[10]~q ),
	.prn(vcc));
defparam \counter[10] .is_wysiwyg = "true";
defparam \counter[10] .power_up = "low";

fiftyfivenm_lcell_comb \Add0~22 (
	.dataa(\counter[11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~21 ),
	.combout(\Add0~22_combout ),
	.cout(\Add0~23 ));
defparam \Add0~22 .lut_mask = 16'h5A5F;
defparam \Add0~22 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \counter[11]~4 (
	.dataa(\Add0~22_combout ),
	.datab(\counter~24_combout ),
	.datac(gnd),
	.datad(\state.GET_WRITE_DATA~q ),
	.cin(gnd),
	.combout(\counter[11]~4_combout ),
	.cout());
defparam \counter[11]~4 .lut_mask = 16'hAACC;
defparam \counter[11]~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add3~22 (
	.dataa(\counter[11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~21 ),
	.combout(\Add3~22_combout ),
	.cout(\Add3~23 ));
defparam \Add3~22 .lut_mask = 16'h5A5F;
defparam \Add3~22 .sum_lutc_input = "cin";

dffeas \counter[11] (
	.clk(clk),
	.d(\counter[11]~4_combout ),
	.asdata(\Add3~22_combout ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.READ_SEND_WAIT~q ),
	.ena(\counter[9]~18_combout ),
	.q(\counter[11]~q ),
	.prn(vcc));
defparam \counter[11] .is_wysiwyg = "true";
defparam \counter[11] .power_up = "low";

fiftyfivenm_lcell_comb \Add0~24 (
	.dataa(\counter[12]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~23 ),
	.combout(\Add0~24_combout ),
	.cout(\Add0~25 ));
defparam \Add0~24 .lut_mask = 16'h5AAF;
defparam \Add0~24 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \counter[12]~3 (
	.dataa(\Add0~24_combout ),
	.datab(\counter~23_combout ),
	.datac(gnd),
	.datad(\state.GET_WRITE_DATA~q ),
	.cin(gnd),
	.combout(\counter[12]~3_combout ),
	.cout());
defparam \counter[12]~3 .lut_mask = 16'hAACC;
defparam \counter[12]~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add3~24 (
	.dataa(\counter[12]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~23 ),
	.combout(\Add3~24_combout ),
	.cout(\Add3~25 ));
defparam \Add3~24 .lut_mask = 16'h5AAF;
defparam \Add3~24 .sum_lutc_input = "cin";

dffeas \counter[12] (
	.clk(clk),
	.d(\counter[12]~3_combout ),
	.asdata(\Add3~24_combout ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.READ_SEND_WAIT~q ),
	.ena(\counter[9]~18_combout ),
	.q(\counter[12]~q ),
	.prn(vcc));
defparam \counter[12] .is_wysiwyg = "true";
defparam \counter[12] .power_up = "low";

fiftyfivenm_lcell_comb \Add0~26 (
	.dataa(\counter[13]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~25 ),
	.combout(\Add0~26_combout ),
	.cout(\Add0~27 ));
defparam \Add0~26 .lut_mask = 16'h5A5F;
defparam \Add0~26 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \counter[13]~2 (
	.dataa(\Add0~26_combout ),
	.datab(\counter~22_combout ),
	.datac(gnd),
	.datad(\state.GET_WRITE_DATA~q ),
	.cin(gnd),
	.combout(\counter[13]~2_combout ),
	.cout());
defparam \counter[13]~2 .lut_mask = 16'hAACC;
defparam \counter[13]~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add3~26 (
	.dataa(\counter[13]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~25 ),
	.combout(\Add3~26_combout ),
	.cout(\Add3~27 ));
defparam \Add3~26 .lut_mask = 16'h5A5F;
defparam \Add3~26 .sum_lutc_input = "cin";

dffeas \counter[13] (
	.clk(clk),
	.d(\counter[13]~2_combout ),
	.asdata(\Add3~26_combout ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.READ_SEND_WAIT~q ),
	.ena(\counter[9]~18_combout ),
	.q(\counter[13]~q ),
	.prn(vcc));
defparam \counter[13] .is_wysiwyg = "true";
defparam \counter[13] .power_up = "low";

fiftyfivenm_lcell_comb \Add0~28 (
	.dataa(\counter[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~27 ),
	.combout(\Add0~28_combout ),
	.cout(\Add0~29 ));
defparam \Add0~28 .lut_mask = 16'h5AAF;
defparam \Add0~28 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \counter[14]~1 (
	.dataa(\Add0~28_combout ),
	.datab(\counter~21_combout ),
	.datac(gnd),
	.datad(\state.GET_WRITE_DATA~q ),
	.cin(gnd),
	.combout(\counter[14]~1_combout ),
	.cout());
defparam \counter[14]~1 .lut_mask = 16'hAACC;
defparam \counter[14]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add3~28 (
	.dataa(\counter[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~27 ),
	.combout(\Add3~28_combout ),
	.cout(\Add3~29 ));
defparam \Add3~28 .lut_mask = 16'h5AAF;
defparam \Add3~28 .sum_lutc_input = "cin";

dffeas \counter[14] (
	.clk(clk),
	.d(\counter[14]~1_combout ),
	.asdata(\Add3~28_combout ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.READ_SEND_WAIT~q ),
	.ena(\counter[9]~18_combout ),
	.q(\counter[14]~q ),
	.prn(vcc));
defparam \counter[14] .is_wysiwyg = "true";
defparam \counter[14] .power_up = "low";

fiftyfivenm_lcell_comb \Add0~30 (
	.dataa(\counter[15]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add0~29 ),
	.combout(\Add0~30_combout ),
	.cout());
defparam \Add0~30 .lut_mask = 16'h5A5A;
defparam \Add0~30 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \counter[15]~0 (
	.dataa(\Add0~30_combout ),
	.datab(\counter~20_combout ),
	.datac(gnd),
	.datad(\state.GET_WRITE_DATA~q ),
	.cin(gnd),
	.combout(\counter[15]~0_combout ),
	.cout());
defparam \counter[15]~0 .lut_mask = 16'hAACC;
defparam \counter[15]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add3~30 (
	.dataa(\counter[15]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add3~29 ),
	.combout(\Add3~30_combout ),
	.cout());
defparam \Add3~30 .lut_mask = 16'h5A5A;
defparam \Add3~30 .sum_lutc_input = "cin";

dffeas \counter[15] (
	.clk(clk),
	.d(\counter[15]~0_combout ),
	.asdata(\Add3~30_combout ),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(\state.READ_SEND_WAIT~q ),
	.ena(\counter[9]~18_combout ),
	.q(\counter[15]~q ),
	.prn(vcc));
defparam \counter[15] .is_wysiwyg = "true";
defparam \counter[15] .power_up = "low";

fiftyfivenm_lcell_comb \Equal10~0 (
	.dataa(\counter[15]~q ),
	.datab(\counter[14]~q ),
	.datac(\counter[13]~q ),
	.datad(\counter[12]~q ),
	.cin(gnd),
	.combout(\Equal10~0_combout ),
	.cout());
defparam \Equal10~0 .lut_mask = 16'h7FFF;
defparam \Equal10~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Equal10~1 (
	.dataa(\counter[8]~q ),
	.datab(\counter[11]~q ),
	.datac(\counter[10]~q ),
	.datad(\counter[9]~q ),
	.cin(gnd),
	.combout(\Equal10~1_combout ),
	.cout());
defparam \Equal10~1 .lut_mask = 16'h7FFF;
defparam \Equal10~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Equal10~2 (
	.dataa(\counter[7]~q ),
	.datab(\counter[6]~q ),
	.datac(\counter[5]~q ),
	.datad(\counter[4]~q ),
	.cin(gnd),
	.combout(\Equal10~2_combout ),
	.cout());
defparam \Equal10~2 .lut_mask = 16'h7FFF;
defparam \Equal10~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Equal10~3 (
	.dataa(\counter[0]~q ),
	.datab(\counter[3]~q ),
	.datac(\counter[2]~q ),
	.datad(\counter[1]~q ),
	.cin(gnd),
	.combout(\Equal10~3_combout ),
	.cout());
defparam \Equal10~3 .lut_mask = 16'hBFFF;
defparam \Equal10~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Equal10~4 (
	.dataa(\Equal10~0_combout ),
	.datab(\Equal10~1_combout ),
	.datac(\Equal10~2_combout ),
	.datad(\Equal10~3_combout ),
	.cin(gnd),
	.combout(\Equal10~4_combout ),
	.cout());
defparam \Equal10~4 .lut_mask = 16'hFFFE;
defparam \Equal10~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \state~68 (
	.dataa(\state.RETURN_PACKET~q ),
	.datab(\Equal10~4_combout ),
	.datac(\state.READ_SEND_WAIT~q ),
	.datad(\out_data[0]~7_combout ),
	.cin(gnd),
	.combout(\state~68_combout ),
	.cout());
defparam \state~68 .lut_mask = 16'hFFFE;
defparam \state~68 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \state~69 (
	.dataa(in_ready),
	.datab(\state~68_combout ),
	.datac(\state.0000~q ),
	.datad(\always1~0_combout ),
	.cin(gnd),
	.combout(\state~69_combout ),
	.cout());
defparam \state~69 .lut_mask = 16'hFFF7;
defparam \state~69 .sum_lutc_input = "datac";

dffeas \state.0000 (
	.clk(clk),
	.d(\state~69_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.0000~q ),
	.prn(vcc));
defparam \state.0000 .is_wysiwyg = "true";
defparam \state.0000 .power_up = "low";

fiftyfivenm_lcell_comb \state~48 (
	.dataa(\state.0000~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\state.GET_WRITE_DATA~q ),
	.cin(gnd),
	.combout(\state~48_combout ),
	.cout());
defparam \state~48 .lut_mask = 16'hAAFF;
defparam \state~48 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \state~65 (
	.dataa(\state~52_combout ),
	.datab(\enable~combout ),
	.datac(\state.GET_ADDR4~q ),
	.datad(\in_ready_0~1_combout ),
	.cin(gnd),
	.combout(\state~65_combout ),
	.cout());
defparam \state~65 .lut_mask = 16'hFEFF;
defparam \state~65 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \state~66 (
	.dataa(\state~64_combout ),
	.datab(\state~48_combout ),
	.datac(\state~65_combout ),
	.datad(\state~53_combout ),
	.cin(gnd),
	.combout(\state~66_combout ),
	.cout());
defparam \state~66 .lut_mask = 16'hFEFF;
defparam \state~66 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \state.GET_EXTRA~2 (
	.dataa(\enable~combout ),
	.datab(out_startofpacket2),
	.datac(\state.GET_EXTRA~q ),
	.datad(\state~66_combout ),
	.cin(gnd),
	.combout(\state.GET_EXTRA~2_combout ),
	.cout());
defparam \state.GET_EXTRA~2 .lut_mask = 16'hFEFF;
defparam \state.GET_EXTRA~2 .sum_lutc_input = "datac";

dffeas \state.GET_EXTRA (
	.clk(clk),
	.d(\state.GET_EXTRA~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.GET_EXTRA~q ),
	.prn(vcc));
defparam \state.GET_EXTRA .is_wysiwyg = "true";
defparam \state.GET_EXTRA .power_up = "low";

fiftyfivenm_lcell_comb \state~73 (
	.dataa(\state.GET_SIZE1~q ),
	.datab(\state.GET_EXTRA~q ),
	.datac(\enable~combout ),
	.datad(out_startofpacket2),
	.cin(gnd),
	.combout(\state~73_combout ),
	.cout());
defparam \state~73 .lut_mask = 16'hACFF;
defparam \state~73 .sum_lutc_input = "datac";

dffeas \state.GET_SIZE1 (
	.clk(clk),
	.d(\state~73_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.GET_SIZE1~q ),
	.prn(vcc));
defparam \state.GET_SIZE1 .is_wysiwyg = "true";
defparam \state.GET_SIZE1 .power_up = "low";

fiftyfivenm_lcell_comb \state~74 (
	.dataa(\state.GET_SIZE2~q ),
	.datab(\state.GET_SIZE1~q ),
	.datac(\enable~combout ),
	.datad(out_startofpacket2),
	.cin(gnd),
	.combout(\state~74_combout ),
	.cout());
defparam \state~74 .lut_mask = 16'hACFF;
defparam \state~74 .sum_lutc_input = "datac";

dffeas \state.GET_SIZE2 (
	.clk(clk),
	.d(\state~74_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.GET_SIZE2~q ),
	.prn(vcc));
defparam \state.GET_SIZE2 .is_wysiwyg = "true";
defparam \state.GET_SIZE2 .power_up = "low";

fiftyfivenm_lcell_comb \state~75 (
	.dataa(\state.GET_ADDR1~q ),
	.datab(\state.GET_SIZE2~q ),
	.datac(\enable~combout ),
	.datad(out_startofpacket2),
	.cin(gnd),
	.combout(\state~75_combout ),
	.cout());
defparam \state~75 .lut_mask = 16'hACFF;
defparam \state~75 .sum_lutc_input = "datac";

dffeas \state.GET_ADDR1 (
	.clk(clk),
	.d(\state~75_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.GET_ADDR1~q ),
	.prn(vcc));
defparam \state.GET_ADDR1 .is_wysiwyg = "true";
defparam \state.GET_ADDR1 .power_up = "low";

fiftyfivenm_lcell_comb \state~76 (
	.dataa(\state.GET_ADDR2~q ),
	.datab(\state.GET_ADDR1~q ),
	.datac(\enable~combout ),
	.datad(out_startofpacket2),
	.cin(gnd),
	.combout(\state~76_combout ),
	.cout());
defparam \state~76 .lut_mask = 16'hACFF;
defparam \state~76 .sum_lutc_input = "datac";

dffeas \state.GET_ADDR2 (
	.clk(clk),
	.d(\state~76_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.GET_ADDR2~q ),
	.prn(vcc));
defparam \state.GET_ADDR2 .is_wysiwyg = "true";
defparam \state.GET_ADDR2 .power_up = "low";

fiftyfivenm_lcell_comb \state~77 (
	.dataa(\state.GET_ADDR3~q ),
	.datab(\state.GET_ADDR2~q ),
	.datac(\enable~combout ),
	.datad(out_startofpacket2),
	.cin(gnd),
	.combout(\state~77_combout ),
	.cout());
defparam \state~77 .lut_mask = 16'hACFF;
defparam \state~77 .sum_lutc_input = "datac";

dffeas \state.GET_ADDR3 (
	.clk(clk),
	.d(\state~77_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.GET_ADDR3~q ),
	.prn(vcc));
defparam \state.GET_ADDR3 .is_wysiwyg = "true";
defparam \state.GET_ADDR3 .power_up = "low";

fiftyfivenm_lcell_comb \state~63 (
	.dataa(\state.GET_ADDR4~q ),
	.datab(\state.GET_ADDR3~q ),
	.datac(\enable~combout ),
	.datad(out_startofpacket2),
	.cin(gnd),
	.combout(\state~63_combout ),
	.cout());
defparam \state~63 .lut_mask = 16'hACFF;
defparam \state~63 .sum_lutc_input = "datac";

dffeas \state.GET_ADDR4 (
	.clk(clk),
	.d(\state~63_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.GET_ADDR4~q ),
	.prn(vcc));
defparam \state.GET_ADDR4 .is_wysiwyg = "true";
defparam \state.GET_ADDR4 .power_up = "low";

fiftyfivenm_lcell_comb \state~72 (
	.dataa(\state.GET_ADDR4~q ),
	.datab(\Equal2~1_combout ),
	.datac(gnd),
	.datad(\command[4]~q ),
	.cin(gnd),
	.combout(\state~72_combout ),
	.cout());
defparam \state~72 .lut_mask = 16'hEEFF;
defparam \state~72 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector1~0 (
	.dataa(\state.GET_WRITE_DATA~q ),
	.datab(\out_data[0]~7_combout ),
	.datac(out_endofpacket2),
	.datad(\enable~combout ),
	.cin(gnd),
	.combout(\Selector1~0_combout ),
	.cout());
defparam \Selector1~0 .lut_mask = 16'hBFFF;
defparam \Selector1~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \in_ready_0~4 (
	.dataa(\last_trans~q ),
	.datab(av_waitrequest),
	.datac(\state.WRITE_WAIT~q ),
	.datad(\Selector1~0_combout ),
	.cin(gnd),
	.combout(\in_ready_0~4_combout ),
	.cout());
defparam \in_ready_0~4 .lut_mask = 16'hEFFF;
defparam \in_ready_0~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \state~81 (
	.dataa(\enable~combout ),
	.datab(out_startofpacket2),
	.datac(\state~72_combout ),
	.datad(\in_ready_0~4_combout ),
	.cin(gnd),
	.combout(\state~81_combout ),
	.cout());
defparam \state~81 .lut_mask = 16'hB1FF;
defparam \state~81 .sum_lutc_input = "datac";

dffeas \state.GET_WRITE_DATA (
	.clk(clk),
	.d(\state~81_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.GET_WRITE_DATA~q ),
	.prn(vcc));
defparam \state.GET_WRITE_DATA .is_wysiwyg = "true";
defparam \state.GET_WRITE_DATA .power_up = "low";

fiftyfivenm_lcell_comb \state~64 (
	.dataa(\enable~combout ),
	.datab(\state.GET_WRITE_DATA~q ),
	.datac(\out_data[0]~7_combout ),
	.datad(out_endofpacket2),
	.cin(gnd),
	.combout(\state~64_combout ),
	.cout());
defparam \state~64 .lut_mask = 16'hFFFE;
defparam \state~64 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \state~67 (
	.dataa(\state~64_combout ),
	.datab(\state.WRITE_WAIT~q ),
	.datac(\state~66_combout ),
	.datad(\always1~0_combout ),
	.cin(gnd),
	.combout(\state~67_combout ),
	.cout());
defparam \state~67 .lut_mask = 16'hEFFF;
defparam \state~67 .sum_lutc_input = "datac";

dffeas \state.WRITE_WAIT (
	.clk(clk),
	.d(\state~67_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.WRITE_WAIT~q ),
	.prn(vcc));
defparam \state.WRITE_WAIT .is_wysiwyg = "true";
defparam \state.WRITE_WAIT .power_up = "low";

fiftyfivenm_lcell_comb \out_data[0]~5 (
	.dataa(\state.WRITE_WAIT~q ),
	.datab(av_waitrequest),
	.datac(gnd),
	.datad(\last_trans~q ),
	.cin(gnd),
	.combout(\out_data[0]~5_combout ),
	.cout());
defparam \out_data[0]~5 .lut_mask = 16'hEEFF;
defparam \out_data[0]~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \WideOr14~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\state.GET_ADDR4~q ),
	.datad(\state.WRITE_WAIT~q ),
	.cin(gnd),
	.combout(\WideOr14~0_combout ),
	.cout());
defparam \WideOr14~0 .lut_mask = 16'h0FFF;
defparam \WideOr14~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \current_byte[1]~1 (
	.dataa(\WideOr14~0_combout ),
	.datab(\current_byte[1]~0_combout ),
	.datac(in_ready),
	.datad(\state.GET_WRITE_DATA~q ),
	.cin(gnd),
	.combout(\current_byte[1]~1_combout ),
	.cout());
defparam \current_byte[1]~1 .lut_mask = 16'h8BFF;
defparam \current_byte[1]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \current_byte[1]~2 (
	.dataa(\out_data[0]~5_combout ),
	.datab(\current_byte[1]~1_combout ),
	.datac(\state.GET_WRITE_DATA~q ),
	.datad(\enable~combout ),
	.cin(gnd),
	.combout(\current_byte[1]~2_combout ),
	.cout());
defparam \current_byte[1]~2 .lut_mask = 16'hFF7F;
defparam \current_byte[1]~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data[0]~6 (
	.dataa(\state.GET_ADDR4~q ),
	.datab(\Equal2~1_combout ),
	.datac(gnd),
	.datad(\enable~combout ),
	.cin(gnd),
	.combout(\out_data[0]~6_combout ),
	.cout());
defparam \out_data[0]~6 .lut_mask = 16'hEEFF;
defparam \out_data[0]~6 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \current_byte[0]~3 (
	.dataa(in_data[0]),
	.datab(\out_data[0]~6_combout ),
	.datac(\current_byte[0]~q ),
	.datad(\state.GET_ADDR4~q ),
	.cin(gnd),
	.combout(\current_byte[0]~3_combout ),
	.cout());
defparam \current_byte[0]~3 .lut_mask = 16'hEFFF;
defparam \current_byte[0]~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \current_byte[0]~4 (
	.dataa(\current_byte[0]~q ),
	.datab(\current_byte[1]~2_combout ),
	.datac(\current_byte[0]~3_combout ),
	.datad(\state.WRITE_WAIT~q ),
	.cin(gnd),
	.combout(\current_byte[0]~4_combout ),
	.cout());
defparam \current_byte[0]~4 .lut_mask = 16'hB8FF;
defparam \current_byte[0]~4 .sum_lutc_input = "datac";

dffeas \current_byte[0] (
	.clk(clk),
	.d(\current_byte[0]~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\current_byte[0]~q ),
	.prn(vcc));
defparam \current_byte[0] .is_wysiwyg = "true";
defparam \current_byte[0] .power_up = "low";

fiftyfivenm_lcell_comb \Selector70~0 (
	.dataa(gnd),
	.datab(\current_byte[1]~q ),
	.datac(\current_byte[0]~q ),
	.datad(\state.GET_ADDR4~q ),
	.cin(gnd),
	.combout(\Selector70~0_combout ),
	.cout());
defparam \Selector70~0 .lut_mask = 16'h3CFF;
defparam \Selector70~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector70~1 (
	.dataa(\Selector70~0_combout ),
	.datab(in_data[1]),
	.datac(\out_data[0]~6_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector70~1_combout ),
	.cout());
defparam \Selector70~1 .lut_mask = 16'hFEFE;
defparam \Selector70~1 .sum_lutc_input = "datac";

dffeas \current_byte[1] (
	.clk(clk),
	.d(\Selector70~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(\state.WRITE_WAIT~q ),
	.sload(gnd),
	.ena(\current_byte[1]~2_combout ),
	.q(\current_byte[1]~q ),
	.prn(vcc));
defparam \current_byte[1] .is_wysiwyg = "true";
defparam \current_byte[1] .power_up = "low";

fiftyfivenm_lcell_comb \Selector82~0 (
	.dataa(\current_byte[1]~q ),
	.datab(\state.RETURN_PACKET~q ),
	.datac(gnd),
	.datad(\current_byte[0]~q ),
	.cin(gnd),
	.combout(\Selector82~0_combout ),
	.cout());
defparam \Selector82~0 .lut_mask = 16'hEEFF;
defparam \Selector82~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_endofpacket~0 (
	.dataa(out_endofpacket1),
	.datab(\Selector82~0_combout ),
	.datac(gnd),
	.datad(in_ready),
	.cin(gnd),
	.combout(\out_endofpacket~0_combout ),
	.cout());
defparam \out_endofpacket~0 .lut_mask = 16'hAACC;
defparam \out_endofpacket~0 .sum_lutc_input = "datac";

dffeas \read_data_buffer[0] (
	.clk(clk),
	.d(readdata[8]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_data~4_combout ),
	.q(\read_data_buffer[0]~q ),
	.prn(vcc));
defparam \read_data_buffer[0] .is_wysiwyg = "true";
defparam \read_data_buffer[0] .power_up = "low";

fiftyfivenm_lcell_comb \out_data[0]~0 (
	.dataa(\state.READ_CMD_WAIT~q ),
	.datab(\state.READ_DATA_WAIT~q ),
	.datac(\current_byte[1]~q ),
	.datad(\state.RETURN_PACKET~q ),
	.cin(gnd),
	.combout(\out_data[0]~0_combout ),
	.cout());
defparam \out_data[0]~0 .lut_mask = 16'hFFFE;
defparam \out_data[0]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data[0]~1 (
	.dataa(\state.RETURN_PACKET~q ),
	.datab(gnd),
	.datac(\state.READ_CMD_WAIT~q ),
	.datad(\state.READ_DATA_WAIT~q ),
	.cin(gnd),
	.combout(\out_data[0]~1_combout ),
	.cout());
defparam \out_data[0]~1 .lut_mask = 16'hAFFF;
defparam \out_data[0]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector80~0 (
	.dataa(\out_data[0]~0_combout ),
	.datab(\counter[8]~q ),
	.datac(\out_data[0]~1_combout ),
	.datad(\command[0]~q ),
	.cin(gnd),
	.combout(\Selector80~0_combout ),
	.cout());
defparam \Selector80~0 .lut_mask = 16'hFFDE;
defparam \Selector80~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector80~1 (
	.dataa(src_data_0),
	.datab(\out_data[0]~0_combout ),
	.datac(\Selector80~0_combout ),
	.datad(\counter[0]~q ),
	.cin(gnd),
	.combout(\Selector80~1_combout ),
	.cout());
defparam \Selector80~1 .lut_mask = 16'hFFBE;
defparam \Selector80~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data[0]~2 (
	.dataa(\out_data[0]~1_combout ),
	.datab(\state.READ_SEND_ISSUE~q ),
	.datac(\out_data[0]~0_combout ),
	.datad(\current_byte[0]~q ),
	.cin(gnd),
	.combout(\out_data[0]~2_combout ),
	.cout());
defparam \out_data[0]~2 .lut_mask = 16'hBFFF;
defparam \out_data[0]~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data[0]~3 (
	.dataa(\out_data[0]~2_combout ),
	.datab(\current_byte[1]~q ),
	.datac(\state.READ_SEND_ISSUE~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_data[0]~3_combout ),
	.cout());
defparam \out_data[0]~3 .lut_mask = 16'hFEFE;
defparam \out_data[0]~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector80~2 (
	.dataa(\read_data_buffer[0]~q ),
	.datab(\Selector80~1_combout ),
	.datac(\state.READ_SEND_ISSUE~q ),
	.datad(\out_data[0]~3_combout ),
	.cin(gnd),
	.combout(\Selector80~2_combout ),
	.cout());
defparam \Selector80~2 .lut_mask = 16'hACFF;
defparam \Selector80~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \WideOr14~1 (
	.dataa(\out_data~4_combout ),
	.datab(\WideOr14~0_combout ),
	.datac(\state.READ_SEND_ISSUE~q ),
	.datad(\state.RETURN_PACKET~q ),
	.cin(gnd),
	.combout(\WideOr14~1_combout ),
	.cout());
defparam \WideOr14~1 .lut_mask = 16'hDFFF;
defparam \WideOr14~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data[0]~8 (
	.dataa(\state.READ_SEND_ISSUE~q ),
	.datab(gnd),
	.datac(\current_byte[1]~q ),
	.datad(\current_byte[0]~q ),
	.cin(gnd),
	.combout(\out_data[0]~8_combout ),
	.cout());
defparam \out_data[0]~8 .lut_mask = 16'hAFFF;
defparam \out_data[0]~8 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data[0]~9 (
	.dataa(in_ready),
	.datab(\out_data[0]~7_combout ),
	.datac(\state.RETURN_PACKET~q ),
	.datad(\out_data[0]~8_combout ),
	.cin(gnd),
	.combout(\out_data[0]~9_combout ),
	.cout());
defparam \out_data[0]~9 .lut_mask = 16'hBFFF;
defparam \out_data[0]~9 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data[0]~10 (
	.dataa(\WideOr14~1_combout ),
	.datab(\out_data[0]~5_combout ),
	.datac(\out_data[0]~6_combout ),
	.datad(\out_data[0]~9_combout ),
	.cin(gnd),
	.combout(\out_data[0]~10_combout ),
	.cout());
defparam \out_data[0]~10 .lut_mask = 16'hFF7F;
defparam \out_data[0]~10 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector72~0 (
	.dataa(out_startofpacket1),
	.datab(\state.READ_SEND_ISSUE~q ),
	.datac(\WideOr14~0_combout ),
	.datad(in_ready),
	.cin(gnd),
	.combout(\Selector72~0_combout ),
	.cout());
defparam \Selector72~0 .lut_mask = 16'hBFFF;
defparam \Selector72~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector38~0 (
	.dataa(\state.GET_ADDR1~q ),
	.datab(\first_trans~q ),
	.datac(gnd),
	.datad(\state.READ_SEND_ISSUE~q ),
	.cin(gnd),
	.combout(\Selector38~0_combout ),
	.cout());
defparam \Selector38~0 .lut_mask = 16'hEEFF;
defparam \Selector38~0 .sum_lutc_input = "datac";

dffeas first_trans(
	.clk(clk),
	.d(\Selector38~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\first_trans~q ),
	.prn(vcc));
defparam first_trans.is_wysiwyg = "true";
defparam first_trans.power_up = "low";

fiftyfivenm_lcell_comb \Selector72~2 (
	.dataa(av_waitrequest),
	.datab(\state.WRITE_WAIT~q ),
	.datac(\last_trans~q ),
	.datad(\Selector72~1_combout ),
	.cin(gnd),
	.combout(\Selector72~2_combout ),
	.cout());
defparam \Selector72~2 .lut_mask = 16'hBFFF;
defparam \Selector72~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector72~3 (
	.dataa(\Selector72~0_combout ),
	.datab(\state.READ_SEND_ISSUE~q ),
	.datac(\first_trans~q ),
	.datad(\Selector72~2_combout ),
	.cin(gnd),
	.combout(\Selector72~3_combout ),
	.cout());
defparam \Selector72~3 .lut_mask = 16'hFEFF;
defparam \Selector72~3 .sum_lutc_input = "datac";

dffeas \read_data_buffer[2] (
	.clk(clk),
	.d(readdata[10]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_data~4_combout ),
	.q(\read_data_buffer[2]~q ),
	.prn(vcc));
defparam \read_data_buffer[2] .is_wysiwyg = "true";
defparam \read_data_buffer[2] .power_up = "low";

dffeas \command[2] (
	.clk(clk),
	.d(in_data[2]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always1~0_combout ),
	.q(\command[2]~q ),
	.prn(vcc));
defparam \command[2] .is_wysiwyg = "true";
defparam \command[2] .power_up = "low";

fiftyfivenm_lcell_comb \Selector78~0 (
	.dataa(\out_data[0]~0_combout ),
	.datab(\counter[10]~q ),
	.datac(\out_data[0]~1_combout ),
	.datad(\command[2]~q ),
	.cin(gnd),
	.combout(\Selector78~0_combout ),
	.cout());
defparam \Selector78~0 .lut_mask = 16'hFFDE;
defparam \Selector78~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector78~1 (
	.dataa(src_data_2),
	.datab(\out_data[0]~0_combout ),
	.datac(\Selector78~0_combout ),
	.datad(\counter[2]~q ),
	.cin(gnd),
	.combout(\Selector78~1_combout ),
	.cout());
defparam \Selector78~1 .lut_mask = 16'hFFBE;
defparam \Selector78~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector78~2 (
	.dataa(\read_data_buffer[2]~q ),
	.datab(\Selector78~1_combout ),
	.datac(\state.READ_SEND_ISSUE~q ),
	.datad(\out_data[0]~3_combout ),
	.cin(gnd),
	.combout(\Selector78~2_combout ),
	.cout());
defparam \Selector78~2 .lut_mask = 16'hACFF;
defparam \Selector78~2 .sum_lutc_input = "datac";

dffeas \read_data_buffer[1] (
	.clk(clk),
	.d(readdata[9]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_data~4_combout ),
	.q(\read_data_buffer[1]~q ),
	.prn(vcc));
defparam \read_data_buffer[1] .is_wysiwyg = "true";
defparam \read_data_buffer[1] .power_up = "low";

fiftyfivenm_lcell_comb \Selector79~0 (
	.dataa(\out_data[0]~1_combout ),
	.datab(src_data_1),
	.datac(\out_data[0]~0_combout ),
	.datad(\command[1]~q ),
	.cin(gnd),
	.combout(\Selector79~0_combout ),
	.cout());
defparam \Selector79~0 .lut_mask = 16'hFFDE;
defparam \Selector79~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector79~1 (
	.dataa(\counter[9]~q ),
	.datab(\out_data[0]~1_combout ),
	.datac(\Selector79~0_combout ),
	.datad(\counter[1]~q ),
	.cin(gnd),
	.combout(\Selector79~1_combout ),
	.cout());
defparam \Selector79~1 .lut_mask = 16'hFFBE;
defparam \Selector79~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector79~2 (
	.dataa(\read_data_buffer[1]~q ),
	.datab(\Selector79~1_combout ),
	.datac(\state.READ_SEND_ISSUE~q ),
	.datad(\out_data[0]~3_combout ),
	.cin(gnd),
	.combout(\Selector79~2_combout ),
	.cout());
defparam \Selector79~2 .lut_mask = 16'hACFF;
defparam \Selector79~2 .sum_lutc_input = "datac";

dffeas \read_data_buffer[5] (
	.clk(clk),
	.d(readdata[13]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_data~4_combout ),
	.q(\read_data_buffer[5]~q ),
	.prn(vcc));
defparam \read_data_buffer[5] .is_wysiwyg = "true";
defparam \read_data_buffer[5] .power_up = "low";

fiftyfivenm_lcell_comb \Selector75~0 (
	.dataa(\out_data[0]~1_combout ),
	.datab(src_payload),
	.datac(\out_data[0]~0_combout ),
	.datad(\command[5]~q ),
	.cin(gnd),
	.combout(\Selector75~0_combout ),
	.cout());
defparam \Selector75~0 .lut_mask = 16'hFFDE;
defparam \Selector75~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector75~1 (
	.dataa(\counter[13]~q ),
	.datab(\out_data[0]~1_combout ),
	.datac(\Selector75~0_combout ),
	.datad(\counter[5]~q ),
	.cin(gnd),
	.combout(\Selector75~1_combout ),
	.cout());
defparam \Selector75~1 .lut_mask = 16'hFFBE;
defparam \Selector75~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector75~2 (
	.dataa(\read_data_buffer[5]~q ),
	.datab(\Selector75~1_combout ),
	.datac(\state.READ_SEND_ISSUE~q ),
	.datad(\out_data[0]~3_combout ),
	.cin(gnd),
	.combout(\Selector75~2_combout ),
	.cout());
defparam \Selector75~2 .lut_mask = 16'hACFF;
defparam \Selector75~2 .sum_lutc_input = "datac";

dffeas \read_data_buffer[7] (
	.clk(clk),
	.d(readdata[15]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_data~4_combout ),
	.q(\read_data_buffer[7]~q ),
	.prn(vcc));
defparam \read_data_buffer[7] .is_wysiwyg = "true";
defparam \read_data_buffer[7] .power_up = "low";

fiftyfivenm_lcell_comb \Selector73~0 (
	.dataa(\state.READ_SEND_ISSUE~q ),
	.datab(\current_byte[0]~q ),
	.datac(\read_data_buffer[7]~q ),
	.datad(\current_byte[1]~q ),
	.cin(gnd),
	.combout(\Selector73~0_combout ),
	.cout());
defparam \Selector73~0 .lut_mask = 16'hFEFF;
defparam \Selector73~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector73~1 (
	.dataa(\Selector73~0_combout ),
	.datab(read_latency_shift_reg_1),
	.datac(readdata_7),
	.datad(\out_data~4_combout ),
	.cin(gnd),
	.combout(\Selector73~1_combout ),
	.cout());
defparam \Selector73~1 .lut_mask = 16'hFFFE;
defparam \Selector73~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector73~2 (
	.dataa(\counter[15]~q ),
	.datab(\counter[7]~q ),
	.datac(\current_byte[1]~q ),
	.datad(\current_byte[0]~q ),
	.cin(gnd),
	.combout(\Selector73~2_combout ),
	.cout());
defparam \Selector73~2 .lut_mask = 16'hEFFE;
defparam \Selector73~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector73~3 (
	.dataa(\Selector73~1_combout ),
	.datab(\state.RETURN_PACKET~q ),
	.datac(in_ready),
	.datad(\Selector73~2_combout ),
	.cin(gnd),
	.combout(\Selector73~3_combout ),
	.cout());
defparam \Selector73~3 .lut_mask = 16'hFFFE;
defparam \Selector73~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \WideOr14~2 (
	.dataa(gnd),
	.datab(\state.RETURN_PACKET~q ),
	.datac(\state.READ_CMD_WAIT~q ),
	.datad(\state.READ_DATA_WAIT~q ),
	.cin(gnd),
	.combout(\WideOr14~2_combout ),
	.cout());
defparam \WideOr14~2 .lut_mask = 16'h3FFF;
defparam \WideOr14~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector73~4 (
	.dataa(\WideOr14~2_combout ),
	.datab(\state.READ_SEND_ISSUE~q ),
	.datac(\WideOr14~0_combout ),
	.datad(\out_data[0]~9_combout ),
	.cin(gnd),
	.combout(\Selector73~4_combout ),
	.cout());
defparam \Selector73~4 .lut_mask = 16'hBFFF;
defparam \Selector73~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector73~5 (
	.dataa(\Selector73~3_combout ),
	.datab(out_data_7),
	.datac(\Selector73~4_combout ),
	.datad(\Selector72~2_combout ),
	.cin(gnd),
	.combout(\Selector73~5_combout ),
	.cout());
defparam \Selector73~5 .lut_mask = 16'hFEFF;
defparam \Selector73~5 .sum_lutc_input = "datac";

dffeas \read_data_buffer[6] (
	.clk(clk),
	.d(readdata[14]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_data~4_combout ),
	.q(\read_data_buffer[6]~q ),
	.prn(vcc));
defparam \read_data_buffer[6] .is_wysiwyg = "true";
defparam \read_data_buffer[6] .power_up = "low";

fiftyfivenm_lcell_comb \Selector74~0 (
	.dataa(\out_data[0]~0_combout ),
	.datab(\counter[14]~q ),
	.datac(\out_data[0]~1_combout ),
	.datad(\command[6]~q ),
	.cin(gnd),
	.combout(\Selector74~0_combout ),
	.cout());
defparam \Selector74~0 .lut_mask = 16'hFFDE;
defparam \Selector74~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector74~1 (
	.dataa(src_payload1),
	.datab(\out_data[0]~0_combout ),
	.datac(\Selector74~0_combout ),
	.datad(\counter[6]~q ),
	.cin(gnd),
	.combout(\Selector74~1_combout ),
	.cout());
defparam \Selector74~1 .lut_mask = 16'hFFBE;
defparam \Selector74~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector74~2 (
	.dataa(\read_data_buffer[6]~q ),
	.datab(\Selector74~1_combout ),
	.datac(\state.READ_SEND_ISSUE~q ),
	.datad(\out_data[0]~3_combout ),
	.cin(gnd),
	.combout(\Selector74~2_combout ),
	.cout());
defparam \Selector74~2 .lut_mask = 16'hACFF;
defparam \Selector74~2 .sum_lutc_input = "datac";

dffeas \read_data_buffer[4] (
	.clk(clk),
	.d(readdata[12]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_data~4_combout ),
	.q(\read_data_buffer[4]~q ),
	.prn(vcc));
defparam \read_data_buffer[4] .is_wysiwyg = "true";
defparam \read_data_buffer[4] .power_up = "low";

fiftyfivenm_lcell_comb \Selector76~0 (
	.dataa(\out_data[0]~0_combout ),
	.datab(\counter[12]~q ),
	.datac(\out_data[0]~1_combout ),
	.datad(\command[4]~q ),
	.cin(gnd),
	.combout(\Selector76~0_combout ),
	.cout());
defparam \Selector76~0 .lut_mask = 16'hFFDE;
defparam \Selector76~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector76~1 (
	.dataa(src_payload2),
	.datab(\out_data[0]~0_combout ),
	.datac(\Selector76~0_combout ),
	.datad(\counter[4]~q ),
	.cin(gnd),
	.combout(\Selector76~1_combout ),
	.cout());
defparam \Selector76~1 .lut_mask = 16'hFFBE;
defparam \Selector76~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector76~2 (
	.dataa(\read_data_buffer[4]~q ),
	.datab(\Selector76~1_combout ),
	.datac(\state.READ_SEND_ISSUE~q ),
	.datad(\out_data[0]~3_combout ),
	.cin(gnd),
	.combout(\Selector76~2_combout ),
	.cout());
defparam \Selector76~2 .lut_mask = 16'hACFF;
defparam \Selector76~2 .sum_lutc_input = "datac";

dffeas \read_data_buffer[3] (
	.clk(clk),
	.d(readdata[11]),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_data~4_combout ),
	.q(\read_data_buffer[3]~q ),
	.prn(vcc));
defparam \read_data_buffer[3] .is_wysiwyg = "true";
defparam \read_data_buffer[3] .power_up = "low";

fiftyfivenm_lcell_comb \Selector77~0 (
	.dataa(\out_data[0]~1_combout ),
	.datab(src_data_3),
	.datac(\out_data[0]~0_combout ),
	.datad(\command[3]~q ),
	.cin(gnd),
	.combout(\Selector77~0_combout ),
	.cout());
defparam \Selector77~0 .lut_mask = 16'hFFDE;
defparam \Selector77~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector77~1 (
	.dataa(\counter[11]~q ),
	.datab(\out_data[0]~1_combout ),
	.datac(\Selector77~0_combout ),
	.datad(\counter[3]~q ),
	.cin(gnd),
	.combout(\Selector77~1_combout ),
	.cout());
defparam \Selector77~1 .lut_mask = 16'hFFBE;
defparam \Selector77~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector77~2 (
	.dataa(\read_data_buffer[3]~q ),
	.datab(\Selector77~1_combout ),
	.datac(\state.READ_SEND_ISSUE~q ),
	.datad(\out_data[0]~3_combout ),
	.cin(gnd),
	.combout(\Selector77~2_combout ),
	.cout());
defparam \Selector77~2 .lut_mask = 16'hACFF;
defparam \Selector77~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector0~0 (
	.dataa(\state.READ_SEND_ISSUE~q ),
	.datab(\state.RETURN_PACKET~q ),
	.datac(\current_byte[1]~q ),
	.datad(\current_byte[0]~q ),
	.cin(gnd),
	.combout(\Selector0~0_combout ),
	.cout());
defparam \Selector0~0 .lut_mask = 16'hEFFF;
defparam \Selector0~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector0~1 (
	.dataa(out_valid1),
	.datab(\state.0000~q ),
	.datac(\WideOr14~0_combout ),
	.datad(\current_byte[1]~0_combout ),
	.cin(gnd),
	.combout(\Selector0~1_combout ),
	.cout());
defparam \Selector0~1 .lut_mask = 16'hEFFF;
defparam \Selector0~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector0~2 (
	.dataa(\Selector0~0_combout ),
	.datab(\Selector0~1_combout ),
	.datac(in_ready),
	.datad(\Selector72~2_combout ),
	.cin(gnd),
	.combout(\Selector0~2_combout ),
	.cout());
defparam \Selector0~2 .lut_mask = 16'hEFFF;
defparam \Selector0~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add2~0 (
	.dataa(\command[2]~q ),
	.datab(address_2),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add2~0_combout ),
	.cout(\Add2~1 ));
defparam \Add2~0 .lut_mask = 16'h66EE;
defparam \Add2~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add2~2 (
	.dataa(address_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~1 ),
	.combout(\Add2~2_combout ),
	.cout(\Add2~3 ));
defparam \Add2~2 .lut_mask = 16'h5A5F;
defparam \Add2~2 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add2~4 (
	.dataa(address_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~3 ),
	.combout(\Add2~4_combout ),
	.cout(\Add2~5 ));
defparam \Add2~4 .lut_mask = 16'h5AAF;
defparam \Add2~4 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add2~6 (
	.dataa(address_5),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~5 ),
	.combout(\Add2~6_combout ),
	.cout(\Add2~7 ));
defparam \Add2~6 .lut_mask = 16'h5A5F;
defparam \Add2~6 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add2~8 (
	.dataa(address_6),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~7 ),
	.combout(\Add2~8_combout ),
	.cout(\Add2~9 ));
defparam \Add2~8 .lut_mask = 16'h5AAF;
defparam \Add2~8 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add2~10 (
	.dataa(address_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~9 ),
	.combout(\Add2~10_combout ),
	.cout(\Add2~11 ));
defparam \Add2~10 .lut_mask = 16'h5A5F;
defparam \Add2~10 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Selector64~0 (
	.dataa(in_data[7]),
	.datab(\Add2~10_combout ),
	.datac(gnd),
	.datad(\state.GET_ADDR4~q ),
	.cin(gnd),
	.combout(\Selector64~0_combout ),
	.cout());
defparam \Selector64~0 .lut_mask = 16'hAACC;
defparam \Selector64~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \address[9]~3 (
	.dataa(\state.WRITE_WAIT~q ),
	.datab(av_waitrequest),
	.datac(\state.READ_SEND_WAIT~q ),
	.datad(\address[9]~2_combout ),
	.cin(gnd),
	.combout(\address[9]~3_combout ),
	.cout());
defparam \address[9]~3 .lut_mask = 16'hFEFF;
defparam \address[9]~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \address[9]~4 (
	.dataa(\state~79_combout ),
	.datab(\Equal10~4_combout ),
	.datac(\state.READ_SEND_WAIT~q ),
	.datad(\address[9]~3_combout ),
	.cin(gnd),
	.combout(\address[9]~4_combout ),
	.cout());
defparam \address[9]~4 .lut_mask = 16'hBFFF;
defparam \address[9]~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \address[4]~6 (
	.dataa(\state.GET_ADDR4~q ),
	.datab(\state.WRITE_WAIT~q ),
	.datac(\state.READ_SEND_WAIT~q ),
	.datad(\address[9]~4_combout ),
	.cin(gnd),
	.combout(\address[4]~6_combout ),
	.cout());
defparam \address[4]~6 .lut_mask = 16'hFFFE;
defparam \address[4]~6 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector65~0 (
	.dataa(in_data[6]),
	.datab(\Add2~8_combout ),
	.datac(gnd),
	.datad(\state.GET_ADDR4~q ),
	.cin(gnd),
	.combout(\Selector65~0_combout ),
	.cout());
defparam \Selector65~0 .lut_mask = 16'hAACC;
defparam \Selector65~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector66~0 (
	.dataa(\Add2~6_combout ),
	.datab(\state.GET_ADDR4~q ),
	.datac(received_esc),
	.datad(out_payload_5),
	.cin(gnd),
	.combout(\Selector66~0_combout ),
	.cout());
defparam \Selector66~0 .lut_mask = 16'hEBBE;
defparam \Selector66~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector67~0 (
	.dataa(in_data[4]),
	.datab(\Add2~4_combout ),
	.datac(gnd),
	.datad(\state.GET_ADDR4~q ),
	.cin(gnd),
	.combout(\Selector67~0_combout ),
	.cout());
defparam \Selector67~0 .lut_mask = 16'hAACC;
defparam \Selector67~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add2~12 (
	.dataa(address_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~11 ),
	.combout(\Add2~12_combout ),
	.cout(\Add2~13 ));
defparam \Add2~12 .lut_mask = 16'h5AAF;
defparam \Add2~12 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add2~14 (
	.dataa(address_9),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add2~13 ),
	.combout(\Add2~14_combout ),
	.cout());
defparam \Add2~14 .lut_mask = 16'h5A5A;
defparam \Add2~14 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Selector62~0 (
	.dataa(in_data[1]),
	.datab(\Add2~14_combout ),
	.datac(gnd),
	.datad(\state.GET_ADDR3~q ),
	.cin(gnd),
	.combout(\Selector62~0_combout ),
	.cout());
defparam \Selector62~0 .lut_mask = 16'hAACC;
defparam \Selector62~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \address[9]~5 (
	.dataa(\state.WRITE_WAIT~q ),
	.datab(\state.READ_SEND_WAIT~q ),
	.datac(\state.GET_ADDR3~q ),
	.datad(\address[9]~4_combout ),
	.cin(gnd),
	.combout(\address[9]~5_combout ),
	.cout());
defparam \address[9]~5 .lut_mask = 16'hFFFE;
defparam \address[9]~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector68~0 (
	.dataa(in_data[3]),
	.datab(\Add2~2_combout ),
	.datac(gnd),
	.datad(\state.GET_ADDR4~q ),
	.cin(gnd),
	.combout(\Selector68~0_combout ),
	.cout());
defparam \Selector68~0 .lut_mask = 16'hAACC;
defparam \Selector68~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector63~0 (
	.dataa(in_data[0]),
	.datab(\Add2~12_combout ),
	.datac(gnd),
	.datad(\state.GET_ADDR3~q ),
	.cin(gnd),
	.combout(\Selector63~0_combout ),
	.cout());
defparam \Selector63~0 .lut_mask = 16'hAACC;
defparam \Selector63~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector81~0 (
	.dataa(av_waitrequest),
	.datab(write1),
	.datac(\state~64_combout ),
	.datad(\state.WRITE_WAIT~q ),
	.cin(gnd),
	.combout(\Selector81~0_combout ),
	.cout());
defparam \Selector81~0 .lut_mask = 16'hFAFC;
defparam \Selector81~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \in_ready_0~2 (
	.dataa(\state.GET_ADDR4~q ),
	.datab(\Equal2~1_combout ),
	.datac(\command[4]~q ),
	.datad(\enable~combout ),
	.cin(gnd),
	.combout(\in_ready_0~2_combout ),
	.cout());
defparam \in_ready_0~2 .lut_mask = 16'hEFFF;
defparam \in_ready_0~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \in_ready_0~3 (
	.dataa(\state.GET_ADDR2~q ),
	.datab(\state.GET_ADDR3~q ),
	.datac(\state.0000~q ),
	.datad(\in_ready_0~0_combout ),
	.cin(gnd),
	.combout(\in_ready_0~3_combout ),
	.cout());
defparam \in_ready_0~3 .lut_mask = 16'hEFFF;
defparam \in_ready_0~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \in_ready_0~5 (
	.dataa(\always1~0_combout ),
	.datab(\in_ready_0~2_combout ),
	.datac(\in_ready_0~3_combout ),
	.datad(\in_ready_0~4_combout ),
	.cin(gnd),
	.combout(\in_ready_0~5_combout ),
	.cout());
defparam \in_ready_0~5 .lut_mask = 16'hFEFF;
defparam \in_ready_0~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector83~0 (
	.dataa(\state.READ_CMD_WAIT~q ),
	.datab(\state.READ_ASSERT~q ),
	.datac(read1),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector83~0_combout ),
	.cout());
defparam \Selector83~0 .lut_mask = 16'hFEFE;
defparam \Selector83~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector83~1 (
	.dataa(\Selector83~0_combout ),
	.datab(av_waitrequest),
	.datac(WideOr1),
	.datad(\state.READ_CMD_WAIT~q ),
	.cin(gnd),
	.combout(\Selector83~1_combout ),
	.cout());
defparam \Selector83~1 .lut_mask = 16'hEFFF;
defparam \Selector83~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector69~0 (
	.dataa(in_data[2]),
	.datab(\Add2~0_combout ),
	.datac(gnd),
	.datad(\state.GET_ADDR4~q ),
	.cin(gnd),
	.combout(\Selector69~0_combout ),
	.cout());
defparam \Selector69~0 .lut_mask = 16'hAACC;
defparam \Selector69~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \writedata[3]~0 (
	.dataa(\state.GET_WRITE_DATA~q ),
	.datab(gnd),
	.datac(\current_byte[1]~q ),
	.datad(\current_byte[0]~q ),
	.cin(gnd),
	.combout(\writedata[3]~0_combout ),
	.cout());
defparam \writedata[3]~0 .lut_mask = 16'hAFFF;
defparam \writedata[3]~0 .sum_lutc_input = "datac";

endmodule

module ADC_altera_avalon_sc_fifo (
	reset,
	out_payload_3,
	out_payload_6,
	out_payload_5,
	out_payload_4,
	out_payload_7,
	out_payload_1,
	out_payload_2,
	out_valid1,
	in_ready_0,
	out_payload_0,
	src_valid,
	src_data_3,
	src_data_6,
	src_data_5,
	src_data_4,
	src_data_7,
	src_data_1,
	src_data_2,
	src_data_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
output 	out_payload_3;
output 	out_payload_6;
output 	out_payload_5;
output 	out_payload_4;
output 	out_payload_7;
output 	out_payload_1;
output 	out_payload_2;
output 	out_valid1;
input 	in_ready_0;
output 	out_payload_0;
input 	src_valid;
input 	src_data_3;
input 	src_data_6;
input 	src_data_5;
input 	src_data_4;
input 	src_data_7;
input 	src_data_1;
input 	src_data_2;
input 	src_data_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_ptr[0]~0_combout ;
wire \wr_ptr[0]~q ;
wire \Add0~5_combout ;
wire \wr_ptr[1]~q ;
wire \internal_out_ready~combout ;
wire \mem_rd_ptr[0]~0_combout ;
wire \rd_ptr[0]~q ;
wire \mem_rd_ptr[1]~1_combout ;
wire \rd_ptr[1]~q ;
wire \internal_out_valid~0_combout ;
wire \Add0~2_combout ;
wire \wr_ptr[2]~q ;
wire \Add0~3_combout ;
wire \wr_ptr[3]~q ;
wire \mem_rd_ptr[3]~3_combout ;
wire \rd_ptr[3]~q ;
wire \Add1~0_combout ;
wire \internal_out_valid~1_combout ;
wire \Add1~1_combout ;
wire \mem_rd_ptr[4]~4_combout ;
wire \rd_ptr[4]~q ;
wire \Add0~0_combout ;
wire \Add0~1_combout ;
wire \wr_ptr[4]~q ;
wire \Add0~4_combout ;
wire \wr_ptr[5]~q ;
wire \mem_rd_ptr[5]~5_combout ;
wire \rd_ptr[5]~q ;
wire \Equal0~0_combout ;
wire \Equal0~1_combout ;
wire \Equal0~2_combout ;
wire \internal_out_valid~2_combout ;
wire \next_empty~0_combout ;
wire \empty~q ;
wire \internal_out_valid~3_combout ;
wire \internal_out_valid~q ;
wire \read~0_combout ;
wire \mem_rd_ptr[2]~2_combout ;
wire \rd_ptr[2]~q ;
wire \next_full~0_combout ;
wire \next_full~1_combout ;
wire \next_full~2_combout ;
wire \next_full~3_combout ;
wire \next_full~4_combout ;
wire \full~q ;
wire \write~combout ;
wire \mem_rtl_0|auto_generated|ram_block1a3~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a6~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a5~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a4~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a7~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a1~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a2~portbdataout ;
wire \mem_rtl_0|auto_generated|ram_block1a0~portbdataout ;

wire [143:0] \mem_rtl_0|auto_generated|ram_block1a3_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a6_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a5_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a7_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a1_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a2_PORTBDATAOUT_bus ;
wire [143:0] \mem_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus ;

assign \mem_rtl_0|auto_generated|ram_block1a3~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a3_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a6~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a6_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a5~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a5_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a4~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a7~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a7_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a1~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a1_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a2~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a2_PORTBDATAOUT_bus [0];

assign \mem_rtl_0|auto_generated|ram_block1a0~portbdataout  = \mem_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus [0];

dffeas \out_payload[3] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a3~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_3),
	.prn(vcc));
defparam \out_payload[3] .is_wysiwyg = "true";
defparam \out_payload[3] .power_up = "low";

dffeas \out_payload[6] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a6~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_6),
	.prn(vcc));
defparam \out_payload[6] .is_wysiwyg = "true";
defparam \out_payload[6] .power_up = "low";

dffeas \out_payload[5] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a5~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_5),
	.prn(vcc));
defparam \out_payload[5] .is_wysiwyg = "true";
defparam \out_payload[5] .power_up = "low";

dffeas \out_payload[4] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a4~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_4),
	.prn(vcc));
defparam \out_payload[4] .is_wysiwyg = "true";
defparam \out_payload[4] .power_up = "low";

dffeas \out_payload[7] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a7~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_7),
	.prn(vcc));
defparam \out_payload[7] .is_wysiwyg = "true";
defparam \out_payload[7] .power_up = "low";

dffeas \out_payload[1] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a1~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_1),
	.prn(vcc));
defparam \out_payload[1] .is_wysiwyg = "true";
defparam \out_payload[1] .power_up = "low";

dffeas \out_payload[2] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a2~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_2),
	.prn(vcc));
defparam \out_payload[2] .is_wysiwyg = "true";
defparam \out_payload[2] .power_up = "low";

dffeas out_valid(
	.clk(clk),
	.d(\internal_out_valid~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_valid1),
	.prn(vcc));
defparam out_valid.is_wysiwyg = "true";
defparam out_valid.power_up = "low";

dffeas \out_payload[0] (
	.clk(clk),
	.d(\mem_rtl_0|auto_generated|ram_block1a0~portbdataout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\internal_out_ready~combout ),
	.q(out_payload_0),
	.prn(vcc));
defparam \out_payload[0] .is_wysiwyg = "true";
defparam \out_payload[0] .power_up = "low";

fiftyfivenm_lcell_comb \wr_ptr[0]~0 (
	.dataa(\wr_ptr[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\wr_ptr[0]~0_combout ),
	.cout());
defparam \wr_ptr[0]~0 .lut_mask = 16'h5555;
defparam \wr_ptr[0]~0 .sum_lutc_input = "datac";

dffeas \wr_ptr[0] (
	.clk(clk),
	.d(\wr_ptr[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~combout ),
	.q(\wr_ptr[0]~q ),
	.prn(vcc));
defparam \wr_ptr[0] .is_wysiwyg = "true";
defparam \wr_ptr[0] .power_up = "low";

fiftyfivenm_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\wr_ptr[0]~q ),
	.datad(\wr_ptr[1]~q ),
	.cin(gnd),
	.combout(\Add0~5_combout ),
	.cout());
defparam \Add0~5 .lut_mask = 16'h0FF0;
defparam \Add0~5 .sum_lutc_input = "datac";

dffeas \wr_ptr[1] (
	.clk(clk),
	.d(\Add0~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~combout ),
	.q(\wr_ptr[1]~q ),
	.prn(vcc));
defparam \wr_ptr[1] .is_wysiwyg = "true";
defparam \wr_ptr[1] .power_up = "low";

fiftyfivenm_lcell_comb internal_out_ready(
	.dataa(in_ready_0),
	.datab(gnd),
	.datac(gnd),
	.datad(out_valid1),
	.cin(gnd),
	.combout(\internal_out_ready~combout ),
	.cout());
defparam internal_out_ready.lut_mask = 16'hAAFF;
defparam internal_out_ready.sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \mem_rd_ptr[0]~0 (
	.dataa(out_valid1),
	.datab(in_ready_0),
	.datac(\rd_ptr[0]~q ),
	.datad(\internal_out_valid~q ),
	.cin(gnd),
	.combout(\mem_rd_ptr[0]~0_combout ),
	.cout());
defparam \mem_rd_ptr[0]~0 .lut_mask = 16'h6996;
defparam \mem_rd_ptr[0]~0 .sum_lutc_input = "datac";

dffeas \rd_ptr[0] (
	.clk(clk),
	.d(\mem_rd_ptr[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_ptr[0]~q ),
	.prn(vcc));
defparam \rd_ptr[0] .is_wysiwyg = "true";
defparam \rd_ptr[0] .power_up = "low";

fiftyfivenm_lcell_comb \mem_rd_ptr[1]~1 (
	.dataa(\rd_ptr[1]~q ),
	.datab(\internal_out_ready~combout ),
	.datac(\internal_out_valid~q ),
	.datad(\rd_ptr[0]~q ),
	.cin(gnd),
	.combout(\mem_rd_ptr[1]~1_combout ),
	.cout());
defparam \mem_rd_ptr[1]~1 .lut_mask = 16'h6996;
defparam \mem_rd_ptr[1]~1 .sum_lutc_input = "datac";

dffeas \rd_ptr[1] (
	.clk(clk),
	.d(\mem_rd_ptr[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_ptr[1]~q ),
	.prn(vcc));
defparam \rd_ptr[1] .is_wysiwyg = "true";
defparam \rd_ptr[1] .power_up = "low";

fiftyfivenm_lcell_comb \internal_out_valid~0 (
	.dataa(\wr_ptr[1]~q ),
	.datab(\rd_ptr[1]~q ),
	.datac(\wr_ptr[0]~q ),
	.datad(\rd_ptr[0]~q ),
	.cin(gnd),
	.combout(\internal_out_valid~0_combout ),
	.cout());
defparam \internal_out_valid~0 .lut_mask = 16'h6996;
defparam \internal_out_valid~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add0~2 (
	.dataa(gnd),
	.datab(\wr_ptr[2]~q ),
	.datac(\wr_ptr[0]~q ),
	.datad(\wr_ptr[1]~q ),
	.cin(gnd),
	.combout(\Add0~2_combout ),
	.cout());
defparam \Add0~2 .lut_mask = 16'hC33C;
defparam \Add0~2 .sum_lutc_input = "datac";

dffeas \wr_ptr[2] (
	.clk(clk),
	.d(\Add0~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~combout ),
	.q(\wr_ptr[2]~q ),
	.prn(vcc));
defparam \wr_ptr[2] .is_wysiwyg = "true";
defparam \wr_ptr[2] .power_up = "low";

fiftyfivenm_lcell_comb \Add0~3 (
	.dataa(\wr_ptr[3]~q ),
	.datab(\wr_ptr[0]~q ),
	.datac(\wr_ptr[1]~q ),
	.datad(\wr_ptr[2]~q ),
	.cin(gnd),
	.combout(\Add0~3_combout ),
	.cout());
defparam \Add0~3 .lut_mask = 16'h6996;
defparam \Add0~3 .sum_lutc_input = "datac";

dffeas \wr_ptr[3] (
	.clk(clk),
	.d(\Add0~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~combout ),
	.q(\wr_ptr[3]~q ),
	.prn(vcc));
defparam \wr_ptr[3] .is_wysiwyg = "true";
defparam \wr_ptr[3] .power_up = "low";

fiftyfivenm_lcell_comb \mem_rd_ptr[3]~3 (
	.dataa(\Add1~0_combout ),
	.datab(\rd_ptr[3]~q ),
	.datac(\internal_out_ready~combout ),
	.datad(\internal_out_valid~q ),
	.cin(gnd),
	.combout(\mem_rd_ptr[3]~3_combout ),
	.cout());
defparam \mem_rd_ptr[3]~3 .lut_mask = 16'hEFFE;
defparam \mem_rd_ptr[3]~3 .sum_lutc_input = "datac";

dffeas \rd_ptr[3] (
	.clk(clk),
	.d(\mem_rd_ptr[3]~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_ptr[3]~q ),
	.prn(vcc));
defparam \rd_ptr[3] .is_wysiwyg = "true";
defparam \rd_ptr[3] .power_up = "low";

fiftyfivenm_lcell_comb \Add1~0 (
	.dataa(\rd_ptr[3]~q ),
	.datab(\rd_ptr[0]~q ),
	.datac(\rd_ptr[1]~q ),
	.datad(\rd_ptr[2]~q ),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout());
defparam \Add1~0 .lut_mask = 16'h6996;
defparam \Add1~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \internal_out_valid~1 (
	.dataa(\read~0_combout ),
	.datab(\internal_out_valid~0_combout ),
	.datac(\wr_ptr[3]~q ),
	.datad(\Add1~0_combout ),
	.cin(gnd),
	.combout(\internal_out_valid~1_combout ),
	.cout());
defparam \internal_out_valid~1 .lut_mask = 16'hEFFE;
defparam \internal_out_valid~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add1~1 (
	.dataa(\rd_ptr[0]~q ),
	.datab(\rd_ptr[1]~q ),
	.datac(\rd_ptr[2]~q ),
	.datad(\rd_ptr[3]~q ),
	.cin(gnd),
	.combout(\Add1~1_combout ),
	.cout());
defparam \Add1~1 .lut_mask = 16'hFFFE;
defparam \Add1~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \mem_rd_ptr[4]~4 (
	.dataa(\rd_ptr[4]~q ),
	.datab(\internal_out_ready~combout ),
	.datac(\internal_out_valid~q ),
	.datad(\Add1~1_combout ),
	.cin(gnd),
	.combout(\mem_rd_ptr[4]~4_combout ),
	.cout());
defparam \mem_rd_ptr[4]~4 .lut_mask = 16'h6996;
defparam \mem_rd_ptr[4]~4 .sum_lutc_input = "datac";

dffeas \rd_ptr[4] (
	.clk(clk),
	.d(\mem_rd_ptr[4]~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_ptr[4]~q ),
	.prn(vcc));
defparam \rd_ptr[4] .is_wysiwyg = "true";
defparam \rd_ptr[4] .power_up = "low";

fiftyfivenm_lcell_comb \Add0~0 (
	.dataa(\wr_ptr[0]~q ),
	.datab(\wr_ptr[1]~q ),
	.datac(\wr_ptr[2]~q ),
	.datad(\wr_ptr[3]~q ),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout());
defparam \Add0~0 .lut_mask = 16'hFFFE;
defparam \Add0~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\wr_ptr[4]~q ),
	.datad(\Add0~0_combout ),
	.cin(gnd),
	.combout(\Add0~1_combout ),
	.cout());
defparam \Add0~1 .lut_mask = 16'h0FF0;
defparam \Add0~1 .sum_lutc_input = "datac";

dffeas \wr_ptr[4] (
	.clk(clk),
	.d(\Add0~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~combout ),
	.q(\wr_ptr[4]~q ),
	.prn(vcc));
defparam \wr_ptr[4] .is_wysiwyg = "true";
defparam \wr_ptr[4] .power_up = "low";

fiftyfivenm_lcell_comb \Add0~4 (
	.dataa(gnd),
	.datab(\wr_ptr[5]~q ),
	.datac(\wr_ptr[4]~q ),
	.datad(\Add0~0_combout ),
	.cin(gnd),
	.combout(\Add0~4_combout ),
	.cout());
defparam \Add0~4 .lut_mask = 16'hC33C;
defparam \Add0~4 .sum_lutc_input = "datac";

dffeas \wr_ptr[5] (
	.clk(clk),
	.d(\Add0~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write~combout ),
	.q(\wr_ptr[5]~q ),
	.prn(vcc));
defparam \wr_ptr[5] .is_wysiwyg = "true";
defparam \wr_ptr[5] .power_up = "low";

fiftyfivenm_lcell_comb \mem_rd_ptr[5]~5 (
	.dataa(\rd_ptr[5]~q ),
	.datab(\read~0_combout ),
	.datac(\rd_ptr[4]~q ),
	.datad(\Add1~1_combout ),
	.cin(gnd),
	.combout(\mem_rd_ptr[5]~5_combout ),
	.cout());
defparam \mem_rd_ptr[5]~5 .lut_mask = 16'h6996;
defparam \mem_rd_ptr[5]~5 .sum_lutc_input = "datac";

dffeas \rd_ptr[5] (
	.clk(clk),
	.d(\mem_rd_ptr[5]~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_ptr[5]~q ),
	.prn(vcc));
defparam \rd_ptr[5] .is_wysiwyg = "true";
defparam \rd_ptr[5] .power_up = "low";

fiftyfivenm_lcell_comb \Equal0~0 (
	.dataa(\rd_ptr[4]~q ),
	.datab(\Add1~1_combout ),
	.datac(\wr_ptr[5]~q ),
	.datad(\rd_ptr[5]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'h6996;
defparam \Equal0~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Equal0~1 (
	.dataa(\rd_ptr[0]~q ),
	.datab(\rd_ptr[1]~q ),
	.datac(\wr_ptr[2]~q ),
	.datad(\rd_ptr[2]~q ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'h6996;
defparam \Equal0~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Equal0~2 (
	.dataa(\wr_ptr[4]~q ),
	.datab(\rd_ptr[4]~q ),
	.datac(\Add1~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal0~2_combout ),
	.cout());
defparam \Equal0~2 .lut_mask = 16'h9696;
defparam \Equal0~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \internal_out_valid~2 (
	.dataa(\internal_out_valid~1_combout ),
	.datab(\Equal0~0_combout ),
	.datac(\Equal0~1_combout ),
	.datad(\Equal0~2_combout ),
	.cin(gnd),
	.combout(\internal_out_valid~2_combout ),
	.cout());
defparam \internal_out_valid~2 .lut_mask = 16'hBFFF;
defparam \internal_out_valid~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \next_empty~0 (
	.dataa(\internal_out_valid~2_combout ),
	.datab(\read~0_combout ),
	.datac(\write~combout ),
	.datad(\empty~q ),
	.cin(gnd),
	.combout(\next_empty~0_combout ),
	.cout());
defparam \next_empty~0 .lut_mask = 16'hFFF7;
defparam \next_empty~0 .sum_lutc_input = "datac";

dffeas empty(
	.clk(clk),
	.d(\next_empty~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\empty~q ),
	.prn(vcc));
defparam empty.is_wysiwyg = "true";
defparam empty.power_up = "low";

fiftyfivenm_lcell_comb \internal_out_valid~3 (
	.dataa(\internal_out_valid~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\empty~q ),
	.cin(gnd),
	.combout(\internal_out_valid~3_combout ),
	.cout());
defparam \internal_out_valid~3 .lut_mask = 16'hFF55;
defparam \internal_out_valid~3 .sum_lutc_input = "datac";

dffeas internal_out_valid(
	.clk(clk),
	.d(\internal_out_valid~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\internal_out_valid~q ),
	.prn(vcc));
defparam internal_out_valid.is_wysiwyg = "true";
defparam internal_out_valid.power_up = "low";

fiftyfivenm_lcell_comb \read~0 (
	.dataa(\internal_out_valid~q ),
	.datab(in_ready_0),
	.datac(gnd),
	.datad(out_valid1),
	.cin(gnd),
	.combout(\read~0_combout ),
	.cout());
defparam \read~0 .lut_mask = 16'hEEFF;
defparam \read~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \mem_rd_ptr[2]~2 (
	.dataa(\rd_ptr[2]~q ),
	.datab(\read~0_combout ),
	.datac(\rd_ptr[0]~q ),
	.datad(\rd_ptr[1]~q ),
	.cin(gnd),
	.combout(\mem_rd_ptr[2]~2_combout ),
	.cout());
defparam \mem_rd_ptr[2]~2 .lut_mask = 16'h6996;
defparam \mem_rd_ptr[2]~2 .sum_lutc_input = "datac";

dffeas \rd_ptr[2] (
	.clk(clk),
	.d(\mem_rd_ptr[2]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\rd_ptr[2]~q ),
	.prn(vcc));
defparam \rd_ptr[2] .is_wysiwyg = "true";
defparam \rd_ptr[2] .power_up = "low";

fiftyfivenm_lcell_comb \next_full~0 (
	.dataa(\rd_ptr[2]~q ),
	.datab(\rd_ptr[4]~q ),
	.datac(\Add0~1_combout ),
	.datad(\Add0~2_combout ),
	.cin(gnd),
	.combout(\next_full~0_combout ),
	.cout());
defparam \next_full~0 .lut_mask = 16'h6996;
defparam \next_full~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \next_full~1 (
	.dataa(\wr_ptr[1]~q ),
	.datab(\rd_ptr[1]~q ),
	.datac(\rd_ptr[0]~q ),
	.datad(\wr_ptr[0]~q ),
	.cin(gnd),
	.combout(\next_full~1_combout ),
	.cout());
defparam \next_full~1 .lut_mask = 16'h6996;
defparam \next_full~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \next_full~2 (
	.dataa(src_valid),
	.datab(\next_full~1_combout ),
	.datac(\rd_ptr[3]~q ),
	.datad(\Add0~3_combout ),
	.cin(gnd),
	.combout(\next_full~2_combout ),
	.cout());
defparam \next_full~2 .lut_mask = 16'hEFFE;
defparam \next_full~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \next_full~3 (
	.dataa(\next_full~0_combout ),
	.datab(\next_full~2_combout ),
	.datac(\rd_ptr[5]~q ),
	.datad(\Add0~4_combout ),
	.cin(gnd),
	.combout(\next_full~3_combout ),
	.cout());
defparam \next_full~3 .lut_mask = 16'hEFFE;
defparam \next_full~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \next_full~4 (
	.dataa(\full~q ),
	.datab(\next_full~3_combout ),
	.datac(gnd),
	.datad(\read~0_combout ),
	.cin(gnd),
	.combout(\next_full~4_combout ),
	.cout());
defparam \next_full~4 .lut_mask = 16'hEEFF;
defparam \next_full~4 .sum_lutc_input = "datac";

dffeas full(
	.clk(clk),
	.d(\next_full~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\full~q ),
	.prn(vcc));
defparam full.is_wysiwyg = "true";
defparam full.power_up = "low";

fiftyfivenm_lcell_comb write(
	.dataa(src_valid),
	.datab(gnd),
	.datac(gnd),
	.datad(\full~q ),
	.cin(gnd),
	.combout(\write~combout ),
	.cout());
defparam write.lut_mask = 16'hAAFF;
defparam write.sum_lutc_input = "datac";

fiftyfivenm_ram_block \mem_rtl_0|auto_generated|ram_block1a3 (
	.portawe(\write~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_3}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~5_combout ,\mem_rd_ptr[4]~4_combout ,\mem_rd_ptr[3]~3_combout ,\mem_rd_ptr[2]~2_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a3_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a3 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .logical_ram_name = "ADC_AvalonBridge:avalonbridge|altera_avalon_sc_fifo:fifo|altsyncram:mem_rtl_0|altsyncram_m4g1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_first_bit_number = 3;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_logical_ram_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_first_bit_number = 3;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_logical_ram_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a3 .ram_block_type = "auto";

fiftyfivenm_ram_block \mem_rtl_0|auto_generated|ram_block1a6 (
	.portawe(\write~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_6}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~5_combout ,\mem_rd_ptr[4]~4_combout ,\mem_rd_ptr[3]~3_combout ,\mem_rd_ptr[2]~2_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a6_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a6 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .logical_ram_name = "ADC_AvalonBridge:avalonbridge|altera_avalon_sc_fifo:fifo|altsyncram:mem_rtl_0|altsyncram_m4g1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_first_bit_number = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_logical_ram_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_first_bit_number = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_logical_ram_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a6 .ram_block_type = "auto";

fiftyfivenm_ram_block \mem_rtl_0|auto_generated|ram_block1a5 (
	.portawe(\write~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_5}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~5_combout ,\mem_rd_ptr[4]~4_combout ,\mem_rd_ptr[3]~3_combout ,\mem_rd_ptr[2]~2_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a5_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a5 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .logical_ram_name = "ADC_AvalonBridge:avalonbridge|altera_avalon_sc_fifo:fifo|altsyncram:mem_rtl_0|altsyncram_m4g1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_first_bit_number = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_logical_ram_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_first_bit_number = 5;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_logical_ram_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a5 .ram_block_type = "auto";

fiftyfivenm_ram_block \mem_rtl_0|auto_generated|ram_block1a4 (
	.portawe(\write~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_4}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~5_combout ,\mem_rd_ptr[4]~4_combout ,\mem_rd_ptr[3]~3_combout ,\mem_rd_ptr[2]~2_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a4 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .logical_ram_name = "ADC_AvalonBridge:avalonbridge|altera_avalon_sc_fifo:fifo|altsyncram:mem_rtl_0|altsyncram_m4g1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_first_bit_number = 4;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_logical_ram_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_first_bit_number = 4;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_logical_ram_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a4 .ram_block_type = "auto";

fiftyfivenm_ram_block \mem_rtl_0|auto_generated|ram_block1a7 (
	.portawe(\write~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_7}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~5_combout ,\mem_rd_ptr[4]~4_combout ,\mem_rd_ptr[3]~3_combout ,\mem_rd_ptr[2]~2_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a7_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a7 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .logical_ram_name = "ADC_AvalonBridge:avalonbridge|altera_avalon_sc_fifo:fifo|altsyncram:mem_rtl_0|altsyncram_m4g1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_first_bit_number = 7;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_logical_ram_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_first_bit_number = 7;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_logical_ram_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a7 .ram_block_type = "auto";

fiftyfivenm_ram_block \mem_rtl_0|auto_generated|ram_block1a1 (
	.portawe(\write~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_1}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~5_combout ,\mem_rd_ptr[4]~4_combout ,\mem_rd_ptr[3]~3_combout ,\mem_rd_ptr[2]~2_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a1_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a1 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .logical_ram_name = "ADC_AvalonBridge:avalonbridge|altera_avalon_sc_fifo:fifo|altsyncram:mem_rtl_0|altsyncram_m4g1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_first_bit_number = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_logical_ram_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_first_bit_number = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_logical_ram_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a1 .ram_block_type = "auto";

fiftyfivenm_ram_block \mem_rtl_0|auto_generated|ram_block1a2 (
	.portawe(\write~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_2}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~5_combout ,\mem_rd_ptr[4]~4_combout ,\mem_rd_ptr[3]~3_combout ,\mem_rd_ptr[2]~2_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a2_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a2 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .logical_ram_name = "ADC_AvalonBridge:avalonbridge|altera_avalon_sc_fifo:fifo|altsyncram:mem_rtl_0|altsyncram_m4g1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_first_bit_number = 2;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_logical_ram_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_first_bit_number = 2;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_logical_ram_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a2 .ram_block_type = "auto";

fiftyfivenm_ram_block \mem_rtl_0|auto_generated|ram_block1a0 (
	.portawe(\write~combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clk),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,src_data_0}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\wr_ptr[5]~q ,\wr_ptr[4]~q ,\wr_ptr[3]~q ,\wr_ptr[2]~q ,\wr_ptr[1]~q ,\wr_ptr[0]~q }),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mem_rd_ptr[5]~5_combout ,\mem_rd_ptr[4]~4_combout ,\mem_rd_ptr[3]~3_combout ,\mem_rd_ptr[2]~2_combout ,\mem_rd_ptr[1]~1_combout ,\mem_rd_ptr[0]~0_combout }),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(\mem_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus ));
defparam \mem_rtl_0|auto_generated|ram_block1a0 .data_interleave_offset_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .data_interleave_width_in_bits = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .logical_ram_name = "ADC_AvalonBridge:avalonbridge|altera_avalon_sc_fifo:fifo|altsyncram:mem_rtl_0|altsyncram_m4g1:auto_generated|ALTSYNCRAM";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .mixed_port_feed_through_mode = "old";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .operation_mode = "dual_port";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_first_bit_number = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_logical_ram_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_address_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_address_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_address_width = 6;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_data_out_clear = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_data_out_clock = "none";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_data_width = 1;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_first_address = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_first_bit_number = 0;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_last_address = 63;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_logical_ram_depth = 64;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_logical_ram_width = 8;
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .port_b_read_enable_clock = "clock0";
defparam \mem_rtl_0|auto_generated|ram_block1a0 .ram_block_type = "auto";

endmodule

module ADC_altera_avalon_st_bytes_to_packets (
	reset_n,
	received_esc1,
	out_payload_3,
	out_payload_6,
	out_payload_5,
	out_payload_4,
	out_payload_7,
	out_payload_1,
	out_payload_2,
	out_valid,
	out_valid1,
	in_ready_0,
	enable,
	out_channel_0,
	out_channel_7,
	out_channel_6,
	out_channel_5,
	out_channel_4,
	out_channel_3,
	out_channel_2,
	out_channel_1,
	received_channel1,
	out_startofpacket1,
	out_endofpacket1,
	out_payload_0,
	out_data_5,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	received_esc1;
input 	out_payload_3;
input 	out_payload_6;
input 	out_payload_5;
input 	out_payload_4;
input 	out_payload_7;
input 	out_payload_1;
input 	out_payload_2;
output 	out_valid;
input 	out_valid1;
input 	in_ready_0;
input 	enable;
output 	out_channel_0;
output 	out_channel_7;
output 	out_channel_6;
output 	out_channel_5;
output 	out_channel_4;
output 	out_channel_3;
output 	out_channel_2;
output 	out_channel_1;
output 	received_channel1;
output 	out_startofpacket1;
output 	out_endofpacket1;
input 	out_payload_0;
output 	out_data_5;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Equal0~0_combout ;
wire \Equal2~0_combout ;
wire \received_esc~0_combout ;
wire \Equal0~1_combout ;
wire \out_channel[7]~2_combout ;
wire \received_channel~0_combout ;
wire \received_channel~1_combout ;
wire \out_startofpacket~0_combout ;
wire \out_startofpacket~1_combout ;
wire \out_endofpacket~0_combout ;
wire \out_endofpacket~1_combout ;


dffeas received_esc(
	.clk(clk),
	.d(\received_esc~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(received_esc1),
	.prn(vcc));
defparam received_esc.is_wysiwyg = "true";
defparam received_esc.power_up = "low";

fiftyfivenm_lcell_comb \out_valid~0 (
	.dataa(received_esc1),
	.datab(gnd),
	.datac(\Equal0~1_combout ),
	.datad(\Equal2~0_combout ),
	.cin(gnd),
	.combout(out_valid),
	.cout());
defparam \out_valid~0 .lut_mask = 16'hAFFF;
defparam \out_valid~0 .sum_lutc_input = "datac";

dffeas \out_channel[0] (
	.clk(clk),
	.d(out_payload_0),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_channel[7]~2_combout ),
	.q(out_channel_0),
	.prn(vcc));
defparam \out_channel[0] .is_wysiwyg = "true";
defparam \out_channel[0] .power_up = "low";

dffeas \out_channel[7] (
	.clk(clk),
	.d(out_payload_7),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_channel[7]~2_combout ),
	.q(out_channel_7),
	.prn(vcc));
defparam \out_channel[7] .is_wysiwyg = "true";
defparam \out_channel[7] .power_up = "low";

dffeas \out_channel[6] (
	.clk(clk),
	.d(out_payload_6),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_channel[7]~2_combout ),
	.q(out_channel_6),
	.prn(vcc));
defparam \out_channel[6] .is_wysiwyg = "true";
defparam \out_channel[6] .power_up = "low";

dffeas \out_channel[5] (
	.clk(clk),
	.d(out_data_5),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_channel[7]~2_combout ),
	.q(out_channel_5),
	.prn(vcc));
defparam \out_channel[5] .is_wysiwyg = "true";
defparam \out_channel[5] .power_up = "low";

dffeas \out_channel[4] (
	.clk(clk),
	.d(out_payload_4),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_channel[7]~2_combout ),
	.q(out_channel_4),
	.prn(vcc));
defparam \out_channel[4] .is_wysiwyg = "true";
defparam \out_channel[4] .power_up = "low";

dffeas \out_channel[3] (
	.clk(clk),
	.d(out_payload_3),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_channel[7]~2_combout ),
	.q(out_channel_3),
	.prn(vcc));
defparam \out_channel[3] .is_wysiwyg = "true";
defparam \out_channel[3] .power_up = "low";

dffeas \out_channel[2] (
	.clk(clk),
	.d(out_payload_2),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_channel[7]~2_combout ),
	.q(out_channel_2),
	.prn(vcc));
defparam \out_channel[2] .is_wysiwyg = "true";
defparam \out_channel[2] .power_up = "low";

dffeas \out_channel[1] (
	.clk(clk),
	.d(out_payload_1),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_channel[7]~2_combout ),
	.q(out_channel_1),
	.prn(vcc));
defparam \out_channel[1] .is_wysiwyg = "true";
defparam \out_channel[1] .power_up = "low";

dffeas received_channel(
	.clk(clk),
	.d(\received_channel~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(received_channel1),
	.prn(vcc));
defparam received_channel.is_wysiwyg = "true";
defparam received_channel.power_up = "low";

dffeas out_startofpacket(
	.clk(clk),
	.d(\out_startofpacket~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(out_startofpacket1),
	.prn(vcc));
defparam out_startofpacket.is_wysiwyg = "true";
defparam out_startofpacket.power_up = "low";

dffeas out_endofpacket(
	.clk(clk),
	.d(\out_endofpacket~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(out_endofpacket1),
	.prn(vcc));
defparam out_endofpacket.is_wysiwyg = "true";
defparam out_endofpacket.power_up = "low";

fiftyfivenm_lcell_comb \out_data[5]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(received_esc1),
	.datad(out_payload_5),
	.cin(gnd),
	.combout(out_data_5),
	.cout());
defparam \out_data[5]~0 .lut_mask = 16'h0FF0;
defparam \out_data[5]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Equal0~0 (
	.dataa(out_payload_6),
	.datab(out_payload_5),
	.datac(out_payload_4),
	.datad(out_payload_7),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hFEFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Equal2~0 (
	.dataa(out_payload_3),
	.datab(\Equal0~0_combout ),
	.datac(out_payload_2),
	.datad(out_payload_1),
	.cin(gnd),
	.combout(\Equal2~0_combout ),
	.cout());
defparam \Equal2~0 .lut_mask = 16'hFEFF;
defparam \Equal2~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \received_esc~0 (
	.dataa(out_payload_0),
	.datab(\Equal2~0_combout ),
	.datac(received_esc1),
	.datad(enable),
	.cin(gnd),
	.combout(\received_esc~0_combout ),
	.cout());
defparam \received_esc~0 .lut_mask = 16'hEFFE;
defparam \received_esc~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Equal0~1 (
	.dataa(out_payload_3),
	.datab(\Equal0~0_combout ),
	.datac(out_payload_1),
	.datad(out_payload_2),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'hFEFF;
defparam \Equal0~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_channel[7]~2 (
	.dataa(out_valid1),
	.datab(in_ready_0),
	.datac(received_channel1),
	.datad(out_valid),
	.cin(gnd),
	.combout(\out_channel[7]~2_combout ),
	.cout());
defparam \out_channel[7]~2 .lut_mask = 16'hFFFE;
defparam \out_channel[7]~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \received_channel~0 (
	.dataa(received_channel1),
	.datab(\Equal2~0_combout ),
	.datac(\Equal0~1_combout ),
	.datad(out_payload_0),
	.cin(gnd),
	.combout(\received_channel~0_combout ),
	.cout());
defparam \received_channel~0 .lut_mask = 16'hFEFF;
defparam \received_channel~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \received_channel~1 (
	.dataa(\received_channel~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(received_esc1),
	.cin(gnd),
	.combout(\received_channel~1_combout ),
	.cout());
defparam \received_channel~1 .lut_mask = 16'hAAFF;
defparam \received_channel~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_startofpacket~0 (
	.dataa(out_startofpacket1),
	.datab(\Equal0~1_combout ),
	.datac(received_esc1),
	.datad(out_payload_0),
	.cin(gnd),
	.combout(\out_startofpacket~0_combout ),
	.cout());
defparam \out_startofpacket~0 .lut_mask = 16'hEFFF;
defparam \out_startofpacket~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_startofpacket~1 (
	.dataa(\out_startofpacket~0_combout ),
	.datab(received_channel1),
	.datac(out_valid),
	.datad(enable),
	.cin(gnd),
	.combout(\out_startofpacket~1_combout ),
	.cout());
defparam \out_startofpacket~1 .lut_mask = 16'hEFFF;
defparam \out_startofpacket~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_endofpacket~0 (
	.dataa(out_endofpacket1),
	.datab(out_payload_0),
	.datac(\Equal0~1_combout ),
	.datad(received_esc1),
	.cin(gnd),
	.combout(\out_endofpacket~0_combout ),
	.cout());
defparam \out_endofpacket~0 .lut_mask = 16'hFEFF;
defparam \out_endofpacket~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_endofpacket~1 (
	.dataa(\out_endofpacket~0_combout ),
	.datab(received_channel1),
	.datac(out_valid),
	.datad(enable),
	.cin(gnd),
	.combout(\out_endofpacket~1_combout ),
	.cout());
defparam \out_endofpacket~1 .lut_mask = 16'hEFFF;
defparam \out_endofpacket~1 .sum_lutc_input = "datac";

endmodule

module ADC_altera_avalon_st_jtag_interface (
	tdo,
	altera_reset_synchronizer_int_chain_out,
	out_data_0,
	out_valid,
	in_data_toggle,
	dreg_6,
	out_data_2,
	out_data_1,
	out_data_6,
	out_data_7,
	out_data_5,
	out_data_3,
	out_data_4,
	src_valid,
	src_data_3,
	src_data_6,
	src_data_5,
	src_data_4,
	src_data_7,
	src_data_1,
	src_data_2,
	src_data_0,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	splitter_nodes_receive_0_3,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	irf_reg_0_1,
	irf_reg_1_1,
	irf_reg_2_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	tdo;
input 	altera_reset_synchronizer_int_chain_out;
input 	out_data_0;
input 	out_valid;
output 	in_data_toggle;
output 	dreg_6;
input 	out_data_2;
input 	out_data_1;
input 	out_data_6;
input 	out_data_7;
input 	out_data_5;
input 	out_data_3;
input 	out_data_4;
output 	src_valid;
output 	src_data_3;
output 	src_data_6;
output 	src_data_5;
output 	src_data_4;
output 	src_data_7;
output 	src_data_1;
output 	src_data_2;
output 	src_data_0;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	splitter_nodes_receive_0_3;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \node|sld_virtual_jtag_component|virtual_state_sdr~0_combout ;
wire \node|sld_virtual_jtag_component|virtual_state_cdr~combout ;
wire \node|sld_virtual_jtag_component|virtual_state_udr~combout ;


ADC_altera_jtag_sld_node node(
	.virtual_state_sdr(\node|sld_virtual_jtag_component|virtual_state_sdr~0_combout ),
	.virtual_state_cdr(\node|sld_virtual_jtag_component|virtual_state_cdr~combout ),
	.virtual_state_udr(\node|sld_virtual_jtag_component|virtual_state_udr~combout ),
	.state_4(state_4),
	.splitter_nodes_receive_0_3(splitter_nodes_receive_0_3),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8));

ADC_altera_jtag_dc_streaming \normal.jtag_dc_streaming (
	.virtual_state_sdr(\node|sld_virtual_jtag_component|virtual_state_sdr~0_combout ),
	.tdo(tdo),
	.virtual_state_cdr(\node|sld_virtual_jtag_component|virtual_state_cdr~combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.virtual_state_udr(\node|sld_virtual_jtag_component|virtual_state_udr~combout ),
	.out_data_0(out_data_0),
	.out_valid(out_valid),
	.in_data_toggle(in_data_toggle),
	.dreg_6(dreg_6),
	.out_data_2(out_data_2),
	.out_data_1(out_data_1),
	.out_data_6(out_data_6),
	.out_data_7(out_data_7),
	.out_data_5(out_data_5),
	.out_data_3(out_data_3),
	.out_data_4(out_data_4),
	.src_valid(src_valid),
	.src_data_3(src_data_3),
	.src_data_6(src_data_6),
	.src_data_5(src_data_5),
	.src_data_4(src_data_4),
	.src_data_7(src_data_7),
	.src_data_1(src_data_1),
	.src_data_2(src_data_2),
	.src_data_0(src_data_0),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.splitter_nodes_receive_0_3(splitter_nodes_receive_0_3),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.irf_reg_0_1(irf_reg_0_1),
	.irf_reg_1_1(irf_reg_1_1),
	.irf_reg_2_1(irf_reg_2_1),
	.clk_clk(clk_clk));

endmodule

module ADC_altera_jtag_dc_streaming (
	virtual_state_sdr,
	tdo,
	virtual_state_cdr,
	altera_reset_synchronizer_int_chain_out,
	virtual_state_udr,
	out_data_0,
	out_valid,
	in_data_toggle,
	dreg_6,
	out_data_2,
	out_data_1,
	out_data_6,
	out_data_7,
	out_data_5,
	out_data_3,
	out_data_4,
	src_valid,
	src_data_3,
	src_data_6,
	src_data_5,
	src_data_4,
	src_data_7,
	src_data_1,
	src_data_2,
	src_data_0,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	splitter_nodes_receive_0_3,
	virtual_ir_scan_reg,
	state_3,
	irf_reg_0_1,
	irf_reg_1_1,
	irf_reg_2_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	virtual_state_sdr;
output 	tdo;
input 	virtual_state_cdr;
input 	altera_reset_synchronizer_int_chain_out;
input 	virtual_state_udr;
input 	out_data_0;
input 	out_valid;
output 	in_data_toggle;
output 	dreg_6;
input 	out_data_2;
input 	out_data_1;
input 	out_data_6;
input 	out_data_7;
input 	out_data_5;
input 	out_data_3;
input 	out_data_4;
output 	src_valid;
output 	src_data_3;
output 	src_data_6;
output 	src_data_5;
output 	src_data_4;
output 	src_data_7;
output 	src_data_1;
output 	src_data_2;
output 	src_data_0;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	splitter_nodes_receive_0_3;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sink_crosser|output_stage|data1[0]~q ;
wire \sink_crosser|output_stage|data1[2]~q ;
wire \sink_crosser|output_stage|data1[1]~q ;
wire \sink_crosser|output_stage|data1[6]~q ;
wire \sink_crosser|output_stage|data1[7]~q ;
wire \sink_crosser|output_stage|data1[5]~q ;
wire \sink_crosser|output_stage|data1[3]~q ;
wire \sink_crosser|output_stage|data1[4]~q ;
wire \jtag_streaming|idle_inserter|out_data~2_combout ;
wire \sink_crosser|output_stage|full1~q ;
wire \synchronizer|dreg[1]~q ;
wire \jtag_streaming|idle_inserter_source_ready~q ;
wire \jtag_streaming|idle_inserter|in_ready~0_combout ;
wire \jtag_streaming|idle_remover_sink_data[3]~q ;
wire \jtag_streaming|idle_remover_sink_data[7]~q ;
wire \jtag_streaming|idle_remover_sink_data[6]~q ;
wire \jtag_streaming|idle_remover_sink_data[4]~q ;
wire \jtag_streaming|idle_remover_sink_data[1]~q ;
wire \jtag_streaming|idle_remover_sink_data[0]~q ;
wire \jtag_streaming|idle_remover_sink_data[2]~q ;
wire \jtag_streaming|idle_remover|out_data[5]~0_combout ;
wire \jtag_streaming|idle_remover|out_valid~combout ;


ADC_altera_jtag_src_crosser source_crosser(
	.sink_reset_n(\synchronizer|dreg[1]~q ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.src_valid1(src_valid),
	.src_data_3(src_data_3),
	.src_data_6(src_data_6),
	.src_data_5(src_data_5),
	.src_data_4(src_data_4),
	.src_data_7(src_data_7),
	.src_data_1(src_data_1),
	.src_data_2(src_data_2),
	.src_data_0(src_data_0),
	.sink_data({\jtag_streaming|idle_remover_sink_data[7]~q ,\jtag_streaming|idle_remover_sink_data[6]~q ,\jtag_streaming|idle_remover|out_data[5]~0_combout ,\jtag_streaming|idle_remover_sink_data[4]~q ,\jtag_streaming|idle_remover_sink_data[3]~q ,
\jtag_streaming|idle_remover_sink_data[2]~q ,\jtag_streaming|idle_remover_sink_data[1]~q ,\jtag_streaming|idle_remover_sink_data[0]~q }),
	.sink_valid(\jtag_streaming|idle_remover|out_valid~combout ),
	.sink_clk(altera_internal_jtag),
	.clk_clk(clk_clk));

ADC_altera_avalon_st_clock_crosser sink_crosser(
	.data1_0(\sink_crosser|output_stage|data1[0]~q ),
	.data1_2(\sink_crosser|output_stage|data1[2]~q ),
	.data1_1(\sink_crosser|output_stage|data1[1]~q ),
	.data1_6(\sink_crosser|output_stage|data1[6]~q ),
	.data1_7(\sink_crosser|output_stage|data1[7]~q ),
	.data1_5(\sink_crosser|output_stage|data1[5]~q ),
	.data1_3(\sink_crosser|output_stage|data1[3]~q ),
	.data1_4(\sink_crosser|output_stage|data1[4]~q ),
	.out_data(\jtag_streaming|idle_inserter|out_data~2_combout ),
	.full1(\sink_crosser|output_stage|full1~q ),
	.dreg_1(\synchronizer|dreg[1]~q ),
	.idle_inserter_source_ready(\jtag_streaming|idle_inserter_source_ready~q ),
	.in_ready(\jtag_streaming|idle_inserter|in_ready~0_combout ),
	.in_reset(altera_reset_synchronizer_int_chain_out),
	.in_data({out_data_7,out_data_6,out_data_5,out_data_4,out_data_3,out_data_2,out_data_1,out_data_0}),
	.out_valid(out_valid),
	.in_data_toggle1(in_data_toggle),
	.dreg_6(dreg_6),
	.altera_internal_jtag(altera_internal_jtag),
	.clk_clk(clk_clk));

ADC_altera_jtag_streaming jtag_streaming(
	.virtual_state_sdr(virtual_state_sdr),
	.tdo(tdo),
	.data1_0(\sink_crosser|output_stage|data1[0]~q ),
	.data1_2(\sink_crosser|output_stage|data1[2]~q ),
	.data1_1(\sink_crosser|output_stage|data1[1]~q ),
	.data1_6(\sink_crosser|output_stage|data1[6]~q ),
	.data1_7(\sink_crosser|output_stage|data1[7]~q ),
	.data1_5(\sink_crosser|output_stage|data1[5]~q ),
	.data1_3(\sink_crosser|output_stage|data1[3]~q ),
	.data1_4(\sink_crosser|output_stage|data1[4]~q ),
	.out_data(\jtag_streaming|idle_inserter|out_data~2_combout ),
	.full1(\sink_crosser|output_stage|full1~q ),
	.reset_n(\synchronizer|dreg[1]~q ),
	.idle_inserter_source_ready1(\jtag_streaming|idle_inserter_source_ready~q ),
	.virtual_state_cdr(virtual_state_cdr),
	.sink_ready(\jtag_streaming|idle_inserter|in_ready~0_combout ),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.virtual_state_udr(virtual_state_udr),
	.idle_remover_sink_data_3(\jtag_streaming|idle_remover_sink_data[3]~q ),
	.idle_remover_sink_data_7(\jtag_streaming|idle_remover_sink_data[7]~q ),
	.idle_remover_sink_data_6(\jtag_streaming|idle_remover_sink_data[6]~q ),
	.idle_remover_sink_data_4(\jtag_streaming|idle_remover_sink_data[4]~q ),
	.idle_remover_sink_data_1(\jtag_streaming|idle_remover_sink_data[1]~q ),
	.idle_remover_sink_data_0(\jtag_streaming|idle_remover_sink_data[0]~q ),
	.idle_remover_sink_data_2(\jtag_streaming|idle_remover_sink_data[2]~q ),
	.out_data_5(\jtag_streaming|idle_remover|out_data[5]~0_combout ),
	.out_valid(\jtag_streaming|idle_remover|out_valid~combout ),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.splitter_nodes_receive_0_3(splitter_nodes_receive_0_3),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.irf_reg_0_1(irf_reg_0_1),
	.irf_reg_1_1(irf_reg_1_1),
	.irf_reg_2_1(irf_reg_2_1),
	.clk_clk(clk_clk));

ADC_altera_std_synchronizer_7 synchronizer(
	.dreg_1(\synchronizer|dreg[1]~q ),
	.reset_n(altera_reset_synchronizer_int_chain_out),
	.clk(altera_internal_jtag));

endmodule

module ADC_altera_avalon_st_clock_crosser (
	data1_0,
	data1_2,
	data1_1,
	data1_6,
	data1_7,
	data1_5,
	data1_3,
	data1_4,
	out_data,
	full1,
	dreg_1,
	idle_inserter_source_ready,
	in_ready,
	in_reset,
	in_data,
	out_valid,
	in_data_toggle1,
	dreg_6,
	altera_internal_jtag,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	data1_0;
output 	data1_2;
output 	data1_1;
output 	data1_6;
output 	data1_7;
output 	data1_5;
output 	data1_3;
output 	data1_4;
input 	out_data;
output 	full1;
input 	dreg_1;
input 	idle_inserter_source_ready;
input 	in_ready;
input 	in_reset;
input 	[7:0] in_data;
input 	out_valid;
output 	in_data_toggle1;
output 	dreg_6;
input 	altera_internal_jtag;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \out_data_buffer[0]~q ;
wire \output_stage|full0~q ;
wire \out_data_buffer[2]~q ;
wire \out_data_buffer[1]~q ;
wire \out_data_buffer[6]~q ;
wire \out_data_buffer[7]~q ;
wire \out_data_buffer[5]~q ;
wire \out_data_buffer[3]~q ;
wire \out_data_buffer[4]~q ;
wire \out_data_toggle_flopped~q ;
wire \in_to_out_synchronizer|dreg[1]~q ;
wire \out_valid_internal~combout ;
wire \in_data_buffer[0]~q ;
wire \in_data_buffer[2]~q ;
wire \in_data_buffer[1]~q ;
wire \in_data_buffer[6]~q ;
wire \in_data_buffer[7]~q ;
wire \in_data_buffer[5]~q ;
wire \in_data_buffer[3]~q ;
wire \in_data_buffer[4]~q ;
wire \out_data_toggle_flopped~0_combout ;
wire \take_in_data~combout ;
wire \in_data_toggle~0_combout ;


ADC_altera_avalon_st_pipeline_base output_stage(
	.data1_0(data1_0),
	.data1_2(data1_2),
	.data1_1(data1_1),
	.data1_6(data1_6),
	.data1_7(data1_7),
	.data1_5(data1_5),
	.data1_3(data1_3),
	.data1_4(data1_4),
	.out_data(out_data),
	.full11(full1),
	.in_data({\out_data_buffer[7]~q ,\out_data_buffer[6]~q ,\out_data_buffer[5]~q ,\out_data_buffer[4]~q ,\out_data_buffer[3]~q ,\out_data_buffer[2]~q ,\out_data_buffer[1]~q ,\out_data_buffer[0]~q }),
	.full01(\output_stage|full0~q ),
	.reset(dreg_1),
	.idle_inserter_source_ready(idle_inserter_source_ready),
	.out_valid_internal(\out_valid_internal~combout ),
	.in_ready(in_ready),
	.clk(altera_internal_jtag));

ADC_altera_std_synchronizer_nocut_1 out_to_in_synchronizer(
	.din(\out_data_toggle_flopped~q ),
	.reset_n(in_reset),
	.dreg_6(dreg_6),
	.clk(clk_clk));

ADC_altera_std_synchronizer_nocut in_to_out_synchronizer(
	.reset_n(dreg_1),
	.dreg_1(\in_to_out_synchronizer|dreg[1]~q ),
	.din(in_data_toggle1),
	.clk(altera_internal_jtag));

dffeas \out_data_buffer[0] (
	.clk(altera_internal_jtag),
	.d(\in_data_buffer[0]~q ),
	.asdata(vcc),
	.clrn(dreg_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_data_buffer[0]~q ),
	.prn(vcc));
defparam \out_data_buffer[0] .is_wysiwyg = "true";
defparam \out_data_buffer[0] .power_up = "low";

dffeas \out_data_buffer[2] (
	.clk(altera_internal_jtag),
	.d(\in_data_buffer[2]~q ),
	.asdata(vcc),
	.clrn(dreg_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_data_buffer[2]~q ),
	.prn(vcc));
defparam \out_data_buffer[2] .is_wysiwyg = "true";
defparam \out_data_buffer[2] .power_up = "low";

dffeas \out_data_buffer[1] (
	.clk(altera_internal_jtag),
	.d(\in_data_buffer[1]~q ),
	.asdata(vcc),
	.clrn(dreg_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_data_buffer[1]~q ),
	.prn(vcc));
defparam \out_data_buffer[1] .is_wysiwyg = "true";
defparam \out_data_buffer[1] .power_up = "low";

dffeas \out_data_buffer[6] (
	.clk(altera_internal_jtag),
	.d(\in_data_buffer[6]~q ),
	.asdata(vcc),
	.clrn(dreg_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_data_buffer[6]~q ),
	.prn(vcc));
defparam \out_data_buffer[6] .is_wysiwyg = "true";
defparam \out_data_buffer[6] .power_up = "low";

dffeas \out_data_buffer[7] (
	.clk(altera_internal_jtag),
	.d(\in_data_buffer[7]~q ),
	.asdata(vcc),
	.clrn(dreg_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_data_buffer[7]~q ),
	.prn(vcc));
defparam \out_data_buffer[7] .is_wysiwyg = "true";
defparam \out_data_buffer[7] .power_up = "low";

dffeas \out_data_buffer[5] (
	.clk(altera_internal_jtag),
	.d(\in_data_buffer[5]~q ),
	.asdata(vcc),
	.clrn(dreg_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_data_buffer[5]~q ),
	.prn(vcc));
defparam \out_data_buffer[5] .is_wysiwyg = "true";
defparam \out_data_buffer[5] .power_up = "low";

dffeas \out_data_buffer[3] (
	.clk(altera_internal_jtag),
	.d(\in_data_buffer[3]~q ),
	.asdata(vcc),
	.clrn(dreg_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_data_buffer[3]~q ),
	.prn(vcc));
defparam \out_data_buffer[3] .is_wysiwyg = "true";
defparam \out_data_buffer[3] .power_up = "low";

dffeas \out_data_buffer[4] (
	.clk(altera_internal_jtag),
	.d(\in_data_buffer[4]~q ),
	.asdata(vcc),
	.clrn(dreg_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_data_buffer[4]~q ),
	.prn(vcc));
defparam \out_data_buffer[4] .is_wysiwyg = "true";
defparam \out_data_buffer[4] .power_up = "low";

dffeas out_data_toggle_flopped(
	.clk(altera_internal_jtag),
	.d(\out_data_toggle_flopped~0_combout ),
	.asdata(vcc),
	.clrn(dreg_1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_data_toggle_flopped~q ),
	.prn(vcc));
defparam out_data_toggle_flopped.is_wysiwyg = "true";
defparam out_data_toggle_flopped.power_up = "low";

fiftyfivenm_lcell_comb out_valid_internal(
	.dataa(gnd),
	.datab(gnd),
	.datac(\out_data_toggle_flopped~q ),
	.datad(\in_to_out_synchronizer|dreg[1]~q ),
	.cin(gnd),
	.combout(\out_valid_internal~combout ),
	.cout());
defparam out_valid_internal.lut_mask = 16'h0FF0;
defparam out_valid_internal.sum_lutc_input = "datac";

dffeas \in_data_buffer[0] (
	.clk(clk_clk),
	.d(in_data[0]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[0]~q ),
	.prn(vcc));
defparam \in_data_buffer[0] .is_wysiwyg = "true";
defparam \in_data_buffer[0] .power_up = "low";

dffeas \in_data_buffer[2] (
	.clk(clk_clk),
	.d(in_data[2]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[2]~q ),
	.prn(vcc));
defparam \in_data_buffer[2] .is_wysiwyg = "true";
defparam \in_data_buffer[2] .power_up = "low";

dffeas \in_data_buffer[1] (
	.clk(clk_clk),
	.d(in_data[1]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[1]~q ),
	.prn(vcc));
defparam \in_data_buffer[1] .is_wysiwyg = "true";
defparam \in_data_buffer[1] .power_up = "low";

dffeas \in_data_buffer[6] (
	.clk(clk_clk),
	.d(in_data[6]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[6]~q ),
	.prn(vcc));
defparam \in_data_buffer[6] .is_wysiwyg = "true";
defparam \in_data_buffer[6] .power_up = "low";

dffeas \in_data_buffer[7] (
	.clk(clk_clk),
	.d(in_data[7]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[7]~q ),
	.prn(vcc));
defparam \in_data_buffer[7] .is_wysiwyg = "true";
defparam \in_data_buffer[7] .power_up = "low";

dffeas \in_data_buffer[5] (
	.clk(clk_clk),
	.d(in_data[5]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[5]~q ),
	.prn(vcc));
defparam \in_data_buffer[5] .is_wysiwyg = "true";
defparam \in_data_buffer[5] .power_up = "low";

dffeas \in_data_buffer[3] (
	.clk(clk_clk),
	.d(in_data[3]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[3]~q ),
	.prn(vcc));
defparam \in_data_buffer[3] .is_wysiwyg = "true";
defparam \in_data_buffer[3] .power_up = "low";

dffeas \in_data_buffer[4] (
	.clk(clk_clk),
	.d(in_data[4]),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\take_in_data~combout ),
	.q(\in_data_buffer[4]~q ),
	.prn(vcc));
defparam \in_data_buffer[4] .is_wysiwyg = "true";
defparam \in_data_buffer[4] .power_up = "low";

fiftyfivenm_lcell_comb \out_data_toggle_flopped~0 (
	.dataa(\out_data_toggle_flopped~q ),
	.datab(\in_to_out_synchronizer|dreg[1]~q ),
	.datac(gnd),
	.datad(\output_stage|full0~q ),
	.cin(gnd),
	.combout(\out_data_toggle_flopped~0_combout ),
	.cout());
defparam \out_data_toggle_flopped~0 .lut_mask = 16'hAACC;
defparam \out_data_toggle_flopped~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb take_in_data(
	.dataa(out_valid),
	.datab(in_data_toggle1),
	.datac(dreg_6),
	.datad(gnd),
	.cin(gnd),
	.combout(\take_in_data~combout ),
	.cout());
defparam take_in_data.lut_mask = 16'hBEBE;
defparam take_in_data.sum_lutc_input = "datac";

dffeas in_data_toggle(
	.clk(clk_clk),
	.d(\in_data_toggle~0_combout ),
	.asdata(vcc),
	.clrn(in_reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(in_data_toggle1),
	.prn(vcc));
defparam in_data_toggle.is_wysiwyg = "true";
defparam in_data_toggle.power_up = "low";

fiftyfivenm_lcell_comb \in_data_toggle~0 (
	.dataa(in_data_toggle1),
	.datab(gnd),
	.datac(out_valid),
	.datad(dreg_6),
	.cin(gnd),
	.combout(\in_data_toggle~0_combout ),
	.cout());
defparam \in_data_toggle~0 .lut_mask = 16'hA0AF;
defparam \in_data_toggle~0 .sum_lutc_input = "datac";

endmodule

module ADC_altera_avalon_st_pipeline_base (
	data1_0,
	data1_2,
	data1_1,
	data1_6,
	data1_7,
	data1_5,
	data1_3,
	data1_4,
	out_data,
	full11,
	in_data,
	full01,
	reset,
	idle_inserter_source_ready,
	out_valid_internal,
	in_ready,
	clk)/* synthesis synthesis_greybox=1 */;
output 	data1_0;
output 	data1_2;
output 	data1_1;
output 	data1_6;
output 	data1_7;
output 	data1_5;
output 	data1_3;
output 	data1_4;
input 	out_data;
output 	full11;
input 	[7:0] in_data;
output 	full01;
input 	reset;
input 	idle_inserter_source_ready;
input 	out_valid_internal;
input 	in_ready;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \data0[0]~q ;
wire \data1~0_combout ;
wire \full0~0_combout ;
wire \data0[2]~q ;
wire \data1~1_combout ;
wire \data0[1]~q ;
wire \data1~2_combout ;
wire \data0[6]~q ;
wire \data1~3_combout ;
wire \data0[7]~q ;
wire \data1~4_combout ;
wire \data0[5]~q ;
wire \data1~5_combout ;
wire \data0[3]~q ;
wire \data1~6_combout ;
wire \data0[4]~q ;
wire \data1~7_combout ;
wire \full1~0_combout ;
wire \full0~1_combout ;


dffeas \data1[0] (
	.clk(clk),
	.d(\data1~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\full0~0_combout ),
	.q(data1_0),
	.prn(vcc));
defparam \data1[0] .is_wysiwyg = "true";
defparam \data1[0] .power_up = "low";

dffeas \data1[2] (
	.clk(clk),
	.d(\data1~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\full0~0_combout ),
	.q(data1_2),
	.prn(vcc));
defparam \data1[2] .is_wysiwyg = "true";
defparam \data1[2] .power_up = "low";

dffeas \data1[1] (
	.clk(clk),
	.d(\data1~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\full0~0_combout ),
	.q(data1_1),
	.prn(vcc));
defparam \data1[1] .is_wysiwyg = "true";
defparam \data1[1] .power_up = "low";

dffeas \data1[6] (
	.clk(clk),
	.d(\data1~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\full0~0_combout ),
	.q(data1_6),
	.prn(vcc));
defparam \data1[6] .is_wysiwyg = "true";
defparam \data1[6] .power_up = "low";

dffeas \data1[7] (
	.clk(clk),
	.d(\data1~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\full0~0_combout ),
	.q(data1_7),
	.prn(vcc));
defparam \data1[7] .is_wysiwyg = "true";
defparam \data1[7] .power_up = "low";

dffeas \data1[5] (
	.clk(clk),
	.d(\data1~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\full0~0_combout ),
	.q(data1_5),
	.prn(vcc));
defparam \data1[5] .is_wysiwyg = "true";
defparam \data1[5] .power_up = "low";

dffeas \data1[3] (
	.clk(clk),
	.d(\data1~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\full0~0_combout ),
	.q(data1_3),
	.prn(vcc));
defparam \data1[3] .is_wysiwyg = "true";
defparam \data1[3] .power_up = "low";

dffeas \data1[4] (
	.clk(clk),
	.d(\data1~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\full0~0_combout ),
	.q(data1_4),
	.prn(vcc));
defparam \data1[4] .is_wysiwyg = "true";
defparam \data1[4] .power_up = "low";

dffeas full1(
	.clk(clk),
	.d(\full1~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!full01),
	.q(full11),
	.prn(vcc));
defparam full1.is_wysiwyg = "true";
defparam full1.power_up = "low";

dffeas full0(
	.clk(clk),
	.d(\full0~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(full01),
	.prn(vcc));
defparam full0.is_wysiwyg = "true";
defparam full0.power_up = "low";

dffeas \data0[0] (
	.clk(clk),
	.d(in_data[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!full01),
	.q(\data0[0]~q ),
	.prn(vcc));
defparam \data0[0] .is_wysiwyg = "true";
defparam \data0[0] .power_up = "low";

fiftyfivenm_lcell_comb \data1~0 (
	.dataa(\data0[0]~q ),
	.datab(in_data[0]),
	.datac(gnd),
	.datad(full01),
	.cin(gnd),
	.combout(\data1~0_combout ),
	.cout());
defparam \data1~0 .lut_mask = 16'hAACC;
defparam \data1~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \full0~0 (
	.dataa(full11),
	.datab(out_data),
	.datac(gnd),
	.datad(idle_inserter_source_ready),
	.cin(gnd),
	.combout(\full0~0_combout ),
	.cout());
defparam \full0~0 .lut_mask = 16'hFF77;
defparam \full0~0 .sum_lutc_input = "datac";

dffeas \data0[2] (
	.clk(clk),
	.d(in_data[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!full01),
	.q(\data0[2]~q ),
	.prn(vcc));
defparam \data0[2] .is_wysiwyg = "true";
defparam \data0[2] .power_up = "low";

fiftyfivenm_lcell_comb \data1~1 (
	.dataa(\data0[2]~q ),
	.datab(in_data[2]),
	.datac(gnd),
	.datad(full01),
	.cin(gnd),
	.combout(\data1~1_combout ),
	.cout());
defparam \data1~1 .lut_mask = 16'hAACC;
defparam \data1~1 .sum_lutc_input = "datac";

dffeas \data0[1] (
	.clk(clk),
	.d(in_data[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!full01),
	.q(\data0[1]~q ),
	.prn(vcc));
defparam \data0[1] .is_wysiwyg = "true";
defparam \data0[1] .power_up = "low";

fiftyfivenm_lcell_comb \data1~2 (
	.dataa(\data0[1]~q ),
	.datab(in_data[1]),
	.datac(gnd),
	.datad(full01),
	.cin(gnd),
	.combout(\data1~2_combout ),
	.cout());
defparam \data1~2 .lut_mask = 16'hAACC;
defparam \data1~2 .sum_lutc_input = "datac";

dffeas \data0[6] (
	.clk(clk),
	.d(in_data[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!full01),
	.q(\data0[6]~q ),
	.prn(vcc));
defparam \data0[6] .is_wysiwyg = "true";
defparam \data0[6] .power_up = "low";

fiftyfivenm_lcell_comb \data1~3 (
	.dataa(\data0[6]~q ),
	.datab(in_data[6]),
	.datac(gnd),
	.datad(full01),
	.cin(gnd),
	.combout(\data1~3_combout ),
	.cout());
defparam \data1~3 .lut_mask = 16'hAACC;
defparam \data1~3 .sum_lutc_input = "datac";

dffeas \data0[7] (
	.clk(clk),
	.d(in_data[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!full01),
	.q(\data0[7]~q ),
	.prn(vcc));
defparam \data0[7] .is_wysiwyg = "true";
defparam \data0[7] .power_up = "low";

fiftyfivenm_lcell_comb \data1~4 (
	.dataa(\data0[7]~q ),
	.datab(in_data[7]),
	.datac(gnd),
	.datad(full01),
	.cin(gnd),
	.combout(\data1~4_combout ),
	.cout());
defparam \data1~4 .lut_mask = 16'hAACC;
defparam \data1~4 .sum_lutc_input = "datac";

dffeas \data0[5] (
	.clk(clk),
	.d(in_data[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!full01),
	.q(\data0[5]~q ),
	.prn(vcc));
defparam \data0[5] .is_wysiwyg = "true";
defparam \data0[5] .power_up = "low";

fiftyfivenm_lcell_comb \data1~5 (
	.dataa(\data0[5]~q ),
	.datab(in_data[5]),
	.datac(gnd),
	.datad(full01),
	.cin(gnd),
	.combout(\data1~5_combout ),
	.cout());
defparam \data1~5 .lut_mask = 16'hAACC;
defparam \data1~5 .sum_lutc_input = "datac";

dffeas \data0[3] (
	.clk(clk),
	.d(in_data[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!full01),
	.q(\data0[3]~q ),
	.prn(vcc));
defparam \data0[3] .is_wysiwyg = "true";
defparam \data0[3] .power_up = "low";

fiftyfivenm_lcell_comb \data1~6 (
	.dataa(\data0[3]~q ),
	.datab(in_data[3]),
	.datac(gnd),
	.datad(full01),
	.cin(gnd),
	.combout(\data1~6_combout ),
	.cout());
defparam \data1~6 .lut_mask = 16'hAACC;
defparam \data1~6 .sum_lutc_input = "datac";

dffeas \data0[4] (
	.clk(clk),
	.d(in_data[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!full01),
	.q(\data0[4]~q ),
	.prn(vcc));
defparam \data0[4] .is_wysiwyg = "true";
defparam \data0[4] .power_up = "low";

fiftyfivenm_lcell_comb \data1~7 (
	.dataa(\data0[4]~q ),
	.datab(in_data[4]),
	.datac(gnd),
	.datad(full01),
	.cin(gnd),
	.combout(\data1~7_combout ),
	.cout());
defparam \data1~7 .lut_mask = 16'hAACC;
defparam \data1~7 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \full1~0 (
	.dataa(out_valid_internal),
	.datab(full11),
	.datac(out_data),
	.datad(idle_inserter_source_ready),
	.cin(gnd),
	.combout(\full1~0_combout ),
	.cout());
defparam \full1~0 .lut_mask = 16'hFEFF;
defparam \full1~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \full0~1 (
	.dataa(full01),
	.datab(out_valid_internal),
	.datac(full11),
	.datad(in_ready),
	.cin(gnd),
	.combout(\full0~1_combout ),
	.cout());
defparam \full0~1 .lut_mask = 16'hACFF;
defparam \full0~1 .sum_lutc_input = "datac";

endmodule

module ADC_altera_std_synchronizer_nocut (
	reset_n,
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module ADC_altera_std_synchronizer_nocut_1 (
	din,
	reset_n,
	dreg_6,
	clk)/* synthesis synthesis_greybox=1 */;
input 	din;
input 	reset_n;
output 	dreg_6;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;
wire \dreg[1]~q ;
wire \dreg[2]~q ;
wire \dreg[3]~q ;
wire \dreg[4]~q ;
wire \dreg[5]~q ;


dffeas \dreg[6] (
	.clk(clk),
	.d(\dreg[5]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_6),
	.prn(vcc));
defparam \dreg[6] .is_wysiwyg = "true";
defparam \dreg[6] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[1]~q ),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas \dreg[2] (
	.clk(clk),
	.d(\dreg[1]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[2]~q ),
	.prn(vcc));
defparam \dreg[2] .is_wysiwyg = "true";
defparam \dreg[2] .power_up = "low";

dffeas \dreg[3] (
	.clk(clk),
	.d(\dreg[2]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[3]~q ),
	.prn(vcc));
defparam \dreg[3] .is_wysiwyg = "true";
defparam \dreg[3] .power_up = "low";

dffeas \dreg[4] (
	.clk(clk),
	.d(\dreg[3]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[4]~q ),
	.prn(vcc));
defparam \dreg[4] .is_wysiwyg = "true";
defparam \dreg[4] .power_up = "low";

dffeas \dreg[5] (
	.clk(clk),
	.d(\dreg[4]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[5]~q ),
	.prn(vcc));
defparam \dreg[5] .is_wysiwyg = "true";
defparam \dreg[5] .power_up = "low";

endmodule

module ADC_altera_jtag_src_crosser (
	sink_reset_n,
	altera_reset_synchronizer_int_chain_out,
	src_valid1,
	src_data_3,
	src_data_6,
	src_data_5,
	src_data_4,
	src_data_7,
	src_data_1,
	src_data_2,
	src_data_0,
	sink_data,
	sink_valid,
	sink_clk,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	sink_reset_n;
input 	altera_reset_synchronizer_int_chain_out;
output 	src_valid1;
output 	src_data_3;
output 	src_data_6;
output 	src_data_5;
output 	src_data_4;
output 	src_data_7;
output 	src_data_1;
output 	src_data_2;
output 	src_data_0;
input 	[7:0] sink_data;
input 	sink_valid;
input 	sink_clk;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \crosser|sync_control_signal~0_combout ;
wire \sink_valid_buffer~q ;
wire \sink_data_buffer[3]~q ;
wire \sink_data_buffer[6]~q ;
wire \sink_data_buffer[5]~q ;
wire \sink_data_buffer[4]~q ;
wire \sink_data_buffer[7]~q ;
wire \sink_data_buffer[1]~q ;
wire \sink_data_buffer[2]~q ;
wire \sink_data_buffer[0]~q ;


ADC_altera_jtag_control_signal_crosser crosser(
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.sync_control_signal(\crosser|sync_control_signal~0_combout ),
	.sink_valid_buffer(\sink_valid_buffer~q ),
	.clk_clk(clk_clk));

dffeas sink_valid_buffer(
	.clk(sink_clk),
	.d(sink_valid),
	.asdata(vcc),
	.clrn(sink_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sink_valid_buffer~q ),
	.prn(vcc));
defparam sink_valid_buffer.is_wysiwyg = "true";
defparam sink_valid_buffer.power_up = "low";

dffeas src_valid(
	.clk(clk_clk),
	.d(\crosser|sync_control_signal~0_combout ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(src_valid1),
	.prn(vcc));
defparam src_valid.is_wysiwyg = "true";
defparam src_valid.power_up = "low";

dffeas \src_data[3] (
	.clk(clk_clk),
	.d(\sink_data_buffer[3]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\crosser|sync_control_signal~0_combout ),
	.q(src_data_3),
	.prn(vcc));
defparam \src_data[3] .is_wysiwyg = "true";
defparam \src_data[3] .power_up = "low";

dffeas \src_data[6] (
	.clk(clk_clk),
	.d(\sink_data_buffer[6]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\crosser|sync_control_signal~0_combout ),
	.q(src_data_6),
	.prn(vcc));
defparam \src_data[6] .is_wysiwyg = "true";
defparam \src_data[6] .power_up = "low";

dffeas \src_data[5] (
	.clk(clk_clk),
	.d(\sink_data_buffer[5]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\crosser|sync_control_signal~0_combout ),
	.q(src_data_5),
	.prn(vcc));
defparam \src_data[5] .is_wysiwyg = "true";
defparam \src_data[5] .power_up = "low";

dffeas \src_data[4] (
	.clk(clk_clk),
	.d(\sink_data_buffer[4]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\crosser|sync_control_signal~0_combout ),
	.q(src_data_4),
	.prn(vcc));
defparam \src_data[4] .is_wysiwyg = "true";
defparam \src_data[4] .power_up = "low";

dffeas \src_data[7] (
	.clk(clk_clk),
	.d(\sink_data_buffer[7]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\crosser|sync_control_signal~0_combout ),
	.q(src_data_7),
	.prn(vcc));
defparam \src_data[7] .is_wysiwyg = "true";
defparam \src_data[7] .power_up = "low";

dffeas \src_data[1] (
	.clk(clk_clk),
	.d(\sink_data_buffer[1]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\crosser|sync_control_signal~0_combout ),
	.q(src_data_1),
	.prn(vcc));
defparam \src_data[1] .is_wysiwyg = "true";
defparam \src_data[1] .power_up = "low";

dffeas \src_data[2] (
	.clk(clk_clk),
	.d(\sink_data_buffer[2]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\crosser|sync_control_signal~0_combout ),
	.q(src_data_2),
	.prn(vcc));
defparam \src_data[2] .is_wysiwyg = "true";
defparam \src_data[2] .power_up = "low";

dffeas \src_data[0] (
	.clk(clk_clk),
	.d(\sink_data_buffer[0]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\crosser|sync_control_signal~0_combout ),
	.q(src_data_0),
	.prn(vcc));
defparam \src_data[0] .is_wysiwyg = "true";
defparam \src_data[0] .power_up = "low";

dffeas \sink_data_buffer[3] (
	.clk(sink_clk),
	.d(sink_data[3]),
	.asdata(vcc),
	.clrn(sink_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sink_valid),
	.q(\sink_data_buffer[3]~q ),
	.prn(vcc));
defparam \sink_data_buffer[3] .is_wysiwyg = "true";
defparam \sink_data_buffer[3] .power_up = "low";

dffeas \sink_data_buffer[6] (
	.clk(sink_clk),
	.d(sink_data[6]),
	.asdata(vcc),
	.clrn(sink_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sink_valid),
	.q(\sink_data_buffer[6]~q ),
	.prn(vcc));
defparam \sink_data_buffer[6] .is_wysiwyg = "true";
defparam \sink_data_buffer[6] .power_up = "low";

dffeas \sink_data_buffer[5] (
	.clk(sink_clk),
	.d(sink_data[5]),
	.asdata(vcc),
	.clrn(sink_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sink_valid),
	.q(\sink_data_buffer[5]~q ),
	.prn(vcc));
defparam \sink_data_buffer[5] .is_wysiwyg = "true";
defparam \sink_data_buffer[5] .power_up = "low";

dffeas \sink_data_buffer[4] (
	.clk(sink_clk),
	.d(sink_data[4]),
	.asdata(vcc),
	.clrn(sink_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sink_valid),
	.q(\sink_data_buffer[4]~q ),
	.prn(vcc));
defparam \sink_data_buffer[4] .is_wysiwyg = "true";
defparam \sink_data_buffer[4] .power_up = "low";

dffeas \sink_data_buffer[7] (
	.clk(sink_clk),
	.d(sink_data[7]),
	.asdata(vcc),
	.clrn(sink_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sink_valid),
	.q(\sink_data_buffer[7]~q ),
	.prn(vcc));
defparam \sink_data_buffer[7] .is_wysiwyg = "true";
defparam \sink_data_buffer[7] .power_up = "low";

dffeas \sink_data_buffer[1] (
	.clk(sink_clk),
	.d(sink_data[1]),
	.asdata(vcc),
	.clrn(sink_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sink_valid),
	.q(\sink_data_buffer[1]~q ),
	.prn(vcc));
defparam \sink_data_buffer[1] .is_wysiwyg = "true";
defparam \sink_data_buffer[1] .power_up = "low";

dffeas \sink_data_buffer[2] (
	.clk(sink_clk),
	.d(sink_data[2]),
	.asdata(vcc),
	.clrn(sink_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sink_valid),
	.q(\sink_data_buffer[2]~q ),
	.prn(vcc));
defparam \sink_data_buffer[2] .is_wysiwyg = "true";
defparam \sink_data_buffer[2] .power_up = "low";

dffeas \sink_data_buffer[0] (
	.clk(sink_clk),
	.d(sink_data[0]),
	.asdata(vcc),
	.clrn(sink_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sink_valid),
	.q(\sink_data_buffer[0]~q ),
	.prn(vcc));
defparam \sink_data_buffer[0] .is_wysiwyg = "true";
defparam \sink_data_buffer[0] .power_up = "low";

endmodule

module ADC_altera_jtag_control_signal_crosser (
	altera_reset_synchronizer_int_chain_out,
	sync_control_signal,
	sink_valid_buffer,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_reset_synchronizer_int_chain_out;
output 	sync_control_signal;
input 	sink_valid_buffer;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \synchronizer|dreg[6]~q ;
wire \edge_detector_register~q ;


ADC_altera_std_synchronizer_2 synchronizer(
	.reset_n(altera_reset_synchronizer_int_chain_out),
	.dreg_6(\synchronizer|dreg[6]~q ),
	.din(sink_valid_buffer),
	.clk(clk_clk));

fiftyfivenm_lcell_comb \sync_control_signal~0 (
	.dataa(\synchronizer|dreg[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\edge_detector_register~q ),
	.cin(gnd),
	.combout(sync_control_signal),
	.cout());
defparam \sync_control_signal~0 .lut_mask = 16'hAAFF;
defparam \sync_control_signal~0 .sum_lutc_input = "datac";

dffeas edge_detector_register(
	.clk(clk_clk),
	.d(\synchronizer|dreg[6]~q ),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\edge_detector_register~q ),
	.prn(vcc));
defparam edge_detector_register.is_wysiwyg = "true";
defparam edge_detector_register.power_up = "low";

endmodule

module ADC_altera_std_synchronizer_2 (
	reset_n,
	dreg_6,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
output 	dreg_6;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;
wire \dreg[1]~q ;
wire \dreg[2]~q ;
wire \dreg[3]~q ;
wire \dreg[4]~q ;
wire \dreg[5]~q ;


dffeas \dreg[6] (
	.clk(clk),
	.d(\dreg[5]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_6),
	.prn(vcc));
defparam \dreg[6] .is_wysiwyg = "true";
defparam \dreg[6] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[1]~q ),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas \dreg[2] (
	.clk(clk),
	.d(\dreg[1]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[2]~q ),
	.prn(vcc));
defparam \dreg[2] .is_wysiwyg = "true";
defparam \dreg[2] .power_up = "low";

dffeas \dreg[3] (
	.clk(clk),
	.d(\dreg[2]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[3]~q ),
	.prn(vcc));
defparam \dreg[3] .is_wysiwyg = "true";
defparam \dreg[3] .power_up = "low";

dffeas \dreg[4] (
	.clk(clk),
	.d(\dreg[3]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[4]~q ),
	.prn(vcc));
defparam \dreg[4] .is_wysiwyg = "true";
defparam \dreg[4] .power_up = "low";

dffeas \dreg[5] (
	.clk(clk),
	.d(\dreg[4]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[5]~q ),
	.prn(vcc));
defparam \dreg[5] .is_wysiwyg = "true";
defparam \dreg[5] .power_up = "low";

endmodule

module ADC_altera_jtag_streaming (
	virtual_state_sdr,
	tdo,
	data1_0,
	data1_2,
	data1_1,
	data1_6,
	data1_7,
	data1_5,
	data1_3,
	data1_4,
	out_data,
	full1,
	reset_n,
	idle_inserter_source_ready1,
	virtual_state_cdr,
	sink_ready,
	altera_reset_synchronizer_int_chain_out,
	virtual_state_udr,
	idle_remover_sink_data_3,
	idle_remover_sink_data_7,
	idle_remover_sink_data_6,
	idle_remover_sink_data_4,
	idle_remover_sink_data_1,
	idle_remover_sink_data_0,
	idle_remover_sink_data_2,
	out_data_5,
	out_valid,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	splitter_nodes_receive_0_3,
	virtual_ir_scan_reg,
	state_3,
	irf_reg_0_1,
	irf_reg_1_1,
	irf_reg_2_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	virtual_state_sdr;
output 	tdo;
input 	data1_0;
input 	data1_2;
input 	data1_1;
input 	data1_6;
input 	data1_7;
input 	data1_5;
input 	data1_3;
input 	data1_4;
output 	out_data;
input 	full1;
input 	reset_n;
output 	idle_inserter_source_ready1;
input 	virtual_state_cdr;
output 	sink_ready;
input 	altera_reset_synchronizer_int_chain_out;
input 	virtual_state_udr;
output 	idle_remover_sink_data_3;
output 	idle_remover_sink_data_7;
output 	idle_remover_sink_data_6;
output 	idle_remover_sink_data_4;
output 	idle_remover_sink_data_1;
output 	idle_remover_sink_data_0;
output 	idle_remover_sink_data_2;
output 	out_data_5;
output 	out_valid;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	splitter_nodes_receive_0_3;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \reset_to_sample_synchronizer|dreg[1]~q ;
wire \idle_inserter|out_data~3_combout ;
wire \clock_to_sample_div2_synchronizer|dreg[1]~q ;
wire \clock_sensor_synchronizer|dreg[1]~q ;
wire \clock_to_sample_div2~q ;
wire \clock_sensor~q ;
wire \idle_inserter|out_data~4_combout ;
wire \clock_sense_reset_n_synchronizer|dreg[6]~q ;
wire \clock_sense_reset_n~q ;
wire \idle_remover_sink_valid~q ;
wire \idle_remover_sink_data[5]~q ;
wire \clock_to_sample_div2~0_combout ;
wire \dr_loopback~0_combout ;
wire \dr_info[4]~2_combout ;
wire \dr_control[0]~1_combout ;
wire \dr_control[8]~q ;
wire \dr_control~8_combout ;
wire \dr_control[7]~q ;
wire \dr_control~7_combout ;
wire \dr_control[6]~q ;
wire \dr_control~6_combout ;
wire \dr_control[5]~q ;
wire \dr_control~5_combout ;
wire \dr_control[4]~q ;
wire \dr_control~4_combout ;
wire \dr_control[3]~q ;
wire \dr_control~3_combout ;
wire \dr_control[2]~q ;
wire \dr_control~2_combout ;
wire \dr_control[1]~q ;
wire \dr_control~0_combout ;
wire \dr_control[0]~q ;
wire \tdo~0_combout ;
wire \dr_debug~3_combout ;
wire \Equal14~2_combout ;
wire \dr_debug[2]~q ;
wire \dr_debug~2_combout ;
wire \dr_debug[0]~1_combout ;
wire \dr_debug[1]~q ;
wire \dr_debug~0_combout ;
wire \dr_debug[0]~q ;
wire \dr_loopback~1_combout ;
wire \dr_loopback~2_combout ;
wire \dr_loopback~q ;
wire \read_data_all_valid~0_combout ;
wire \Equal14~0_combout ;
wire \offset[7]~0_combout ;
wire \offset[2]~q ;
wire \offset[1]~q ;
wire \offset[0]~q ;
wire \Equal6~0_combout ;
wire \offset[3]~q ;
wire \offset[4]~q ;
wire \offset[5]~q ;
wire \offset[6]~q ;
wire \Equal6~1_combout ;
wire \offset[7]~q ;
wire \Equal6~2_combout ;
wire \write_state~22_combout ;
wire \write_state~19_combout ;
wire \write_state.ST_BYPASS~q ;
wire \bypass_bit_counter[0]~8_combout ;
wire \bypass_bit_counter~12_combout ;
wire \bypass_bit_counter[0]~13_combout ;
wire \bypass_bit_counter[0]~q ;
wire \bypass_bit_counter[0]~9 ;
wire \bypass_bit_counter[1]~10_combout ;
wire \bypass_bit_counter[1]~q ;
wire \bypass_bit_counter[1]~11 ;
wire \bypass_bit_counter[2]~14_combout ;
wire \bypass_bit_counter[2]~q ;
wire \write_state~14_combout ;
wire \bypass_bit_counter[2]~15 ;
wire \bypass_bit_counter[3]~16_combout ;
wire \bypass_bit_counter[3]~q ;
wire \bypass_bit_counter[3]~17 ;
wire \bypass_bit_counter[4]~18_combout ;
wire \bypass_bit_counter[4]~q ;
wire \bypass_bit_counter[4]~19 ;
wire \bypass_bit_counter[5]~20_combout ;
wire \bypass_bit_counter[5]~q ;
wire \bypass_bit_counter[5]~21 ;
wire \bypass_bit_counter[6]~22_combout ;
wire \bypass_bit_counter[6]~q ;
wire \bypass_bit_counter[6]~23 ;
wire \bypass_bit_counter[7]~24_combout ;
wire \bypass_bit_counter[7]~q ;
wire \write_state~15_combout ;
wire \write_state~16_combout ;
wire \write_state~18_combout ;
wire \write_state.ST_HEADER_2~q ;
wire \write_state~21_combout ;
wire \write_state.ST_WRITE_DATA~q ;
wire \header_in_bit_counter~3_combout ;
wire \header_in_bit_counter[0]~4_combout ;
wire \header_in_bit_counter[0]~5_combout ;
wire \header_in_bit_counter[0]~q ;
wire \header_in_bit_counter~2_combout ;
wire \header_in_bit_counter~6_combout ;
wire \header_in_bit_counter[1]~q ;
wire \header_in_bit_counter~8_combout ;
wire \header_in_bit_counter[2]~q ;
wire \Add1~0_combout ;
wire \header_in_bit_counter~7_combout ;
wire \header_in_bit_counter[3]~q ;
wire \read_data_length[0]~0_combout ;
wire \read_data_length[0]~2_combout ;
wire \write_data_length[0]~0_combout ;
wire \write_state~17_combout ;
wire \write_state~20_combout ;
wire \write_state.ST_HEADER_1~q ;
wire \read_data_length[0]~1_combout ;
wire \read_data_length[2]~q ;
wire \header_in[14]~0_combout ;
wire \header_in[15]~q ;
wire \header_in[14]~q ;
wire \read_data_length[0]~q ;
wire \read_data_length[1]~q ;
wire \read_data_all_valid~1_combout ;
wire \decode_header_1~2_combout ;
wire \decode_header_1~3_combout ;
wire \decode_header_1~q ;
wire \read_data_all_valid~2_combout ;
wire \read_data_all_valid~3_combout ;
wire \read_data_all_valid~q ;
wire \Add8~0_combout ;
wire \header_out_bit_counter~0_combout ;
wire \header_out_bit_counter[0]~1_combout ;
wire \header_out_bit_counter[0]~q ;
wire \header_out_bit_counter~4_combout ;
wire \header_out_bit_counter[1]~q ;
wire \Add6~0_combout ;
wire \header_out_bit_counter~2_combout ;
wire \header_out_bit_counter[2]~q ;
wire \Add6~1_combout ;
wire \header_out_bit_counter~3_combout ;
wire \header_out_bit_counter[3]~q ;
wire \Equal16~0_combout ;
wire \read_state~11_combout ;
wire \read_state~12_combout ;
wire \dr_data_out[2]~18_combout ;
wire \read_state~14_combout ;
wire \read_state~9_combout ;
wire \read_state~10_combout ;
wire \read_state.ST_PADDED~q ;
wire \read_state~8_combout ;
wire \read_state.ST_READ_DATA~q ;
wire \read_state~13_combout ;
wire \read_state.ST_HEADER~q ;
wire \padded_bit_counter[0]~0_combout ;
wire \padded_bit_counter~1_combout ;
wire \padded_bit_counter[0]~2_combout ;
wire \padded_bit_counter[0]~q ;
wire \Add8~1 ;
wire \Add8~2_combout ;
wire \padded_bit_counter~3_combout ;
wire \padded_bit_counter[1]~q ;
wire \Add8~3 ;
wire \Add8~4_combout ;
wire \padded_bit_counter~4_combout ;
wire \padded_bit_counter[2]~q ;
wire \Add5~0_combout ;
wire \Add8~5 ;
wire \Add8~6_combout ;
wire \padded_bit_counter~5_combout ;
wire \padded_bit_counter[3]~q ;
wire \Add5~1 ;
wire \Add5~2_combout ;
wire \Add8~7 ;
wire \Add8~8_combout ;
wire \padded_bit_counter~6_combout ;
wire \padded_bit_counter[4]~q ;
wire \idle_inserter_source_ready~0_combout ;
wire \Add5~3 ;
wire \Add5~4_combout ;
wire \Add8~9 ;
wire \Add8~10_combout ;
wire \padded_bit_counter~7_combout ;
wire \padded_bit_counter[5]~q ;
wire \Add5~5 ;
wire \Add5~6_combout ;
wire \Add8~11 ;
wire \Add8~12_combout ;
wire \padded_bit_counter~8_combout ;
wire \padded_bit_counter[6]~q ;
wire \Add5~7 ;
wire \Add5~8_combout ;
wire \Add8~13 ;
wire \Add8~14_combout ;
wire \padded_bit_counter~9_combout ;
wire \padded_bit_counter[7]~q ;
wire \Add5~9 ;
wire \Add5~10_combout ;
wire \padded_bit_counter~10_combout ;
wire \Add8~15 ;
wire \Add8~16_combout ;
wire \dr_data_out[2]~11_combout ;
wire \padded_bit_counter~11_combout ;
wire \padded_bit_counter[8]~q ;
wire \idle_inserter_source_ready~1_combout ;
wire \Equal17~0_combout ;
wire \dr_data_out~7_combout ;
wire \read_data_bit_counter~0_combout ;
wire \read_data_bit_counter[0]~1_combout ;
wire \read_data_bit_counter[0]~q ;
wire \read_data_bit_counter~2_combout ;
wire \read_data_bit_counter[1]~q ;
wire \Add9~0_combout ;
wire \read_data_bit_counter~3_combout ;
wire \read_data_bit_counter[2]~q ;
wire \Equal1~0_combout ;
wire \dr_data_out[2]~12_combout ;
wire \dr_data_out[2]~13_combout ;
wire \Add10~0_combout ;
wire \scan_length_byte_counter[0]~21_combout ;
wire \scan_length_byte_counter[0]~q ;
wire \Add10~1 ;
wire \Add10~2_combout ;
wire \scan_length_byte_counter[1]~13_combout ;
wire \scan_length_byte_counter[1]~q ;
wire \Add10~3 ;
wire \Add10~4_combout ;
wire \scan_length_byte_counter[2]~14_combout ;
wire \scan_length_byte_counter[2]~q ;
wire \Add10~5 ;
wire \Add10~6_combout ;
wire \scan_length_byte_counter[3]~15_combout ;
wire \scan_length_byte_counter[3]~q ;
wire \Add10~7 ;
wire \Add10~8_combout ;
wire \scan_length_byte_counter[4]~16_combout ;
wire \scan_length_byte_counter[4]~q ;
wire \Equal3~1_combout ;
wire \Add10~9 ;
wire \Add10~10_combout ;
wire \scan_length_byte_counter[5]~17_combout ;
wire \scan_length_byte_counter[5]~q ;
wire \Add10~11 ;
wire \Add10~12_combout ;
wire \scan_length_byte_counter[6]~18_combout ;
wire \scan_length_byte_counter[6]~q ;
wire \Equal3~2_combout ;
wire \Equal3~0_combout ;
wire \Add10~29 ;
wire \Add10~30_combout ;
wire \header_in[13]~q ;
wire \header_in[12]~q ;
wire \header_in[11]~q ;
wire \scan_length[7]~q ;
wire \scan_length_byte_counter[15]~7_combout ;
wire \scan_length_byte_counter[15]~q ;
wire \Add10~31 ;
wire \Add10~32_combout ;
wire \scan_length[8]~q ;
wire \scan_length_byte_counter[16]~8_combout ;
wire \scan_length_byte_counter[16]~q ;
wire \Add10~33 ;
wire \Add10~34_combout ;
wire \scan_length[9]~q ;
wire \scan_length_byte_counter[17]~9_combout ;
wire \scan_length_byte_counter[17]~q ;
wire \Add10~35 ;
wire \Add10~36_combout ;
wire \scan_length_byte_counter[18]~20_combout ;
wire \scan_length_byte_counter[18]~q ;
wire \Equal3~3_combout ;
wire \Equal3~4_combout ;
wire \scan_length_byte_counter[1]~10_combout ;
wire \scan_length_byte_counter[1]~11_combout ;
wire \scan_length_byte_counter[0]~12_combout ;
wire \Add10~13 ;
wire \Add10~14_combout ;
wire \scan_length_byte_counter[7]~19_combout ;
wire \scan_length_byte_counter[7]~q ;
wire \Add10~15 ;
wire \Add10~16_combout ;
wire \header_in[10]~q ;
wire \header_in[9]~q ;
wire \header_in[8]~q ;
wire \header_in[7]~q ;
wire \header_in[6]~q ;
wire \header_in[5]~q ;
wire \header_in[4]~q ;
wire \scan_length[0]~q ;
wire \scan_length_byte_counter[8]~0_combout ;
wire \scan_length_byte_counter[8]~q ;
wire \Add10~17 ;
wire \Add10~18_combout ;
wire \scan_length[1]~q ;
wire \scan_length_byte_counter[9]~1_combout ;
wire \scan_length_byte_counter[9]~q ;
wire \Add10~19 ;
wire \Add10~20_combout ;
wire \scan_length[2]~q ;
wire \scan_length_byte_counter[10]~2_combout ;
wire \scan_length_byte_counter[10]~q ;
wire \Add10~21 ;
wire \Add10~22_combout ;
wire \scan_length[3]~q ;
wire \scan_length_byte_counter[11]~3_combout ;
wire \scan_length_byte_counter[11]~q ;
wire \Add10~23 ;
wire \Add10~24_combout ;
wire \scan_length[4]~q ;
wire \scan_length_byte_counter[12]~4_combout ;
wire \scan_length_byte_counter[12]~q ;
wire \Add10~25 ;
wire \Add10~26_combout ;
wire \scan_length[5]~q ;
wire \scan_length_byte_counter[13]~5_combout ;
wire \scan_length_byte_counter[13]~q ;
wire \Add10~27 ;
wire \Add10~28_combout ;
wire \scan_length[6]~q ;
wire \scan_length_byte_counter[14]~6_combout ;
wire \scan_length_byte_counter[14]~q ;
wire \decoded_read_data_length[13]~0_combout ;
wire \decoded_read_data_length[12]~1_combout ;
wire \decoded_read_data_length[11]~2_combout ;
wire \decoded_read_data_length[10]~3_combout ;
wire \decoded_read_data_length[9]~4_combout ;
wire \decoded_read_data_length[8]~5_combout ;
wire \LessThan0~1_cout ;
wire \LessThan0~3_cout ;
wire \LessThan0~5_cout ;
wire \LessThan0~7_cout ;
wire \LessThan0~9_cout ;
wire \LessThan0~11_cout ;
wire \LessThan0~13_cout ;
wire \LessThan0~14_combout ;
wire \read_data_valid~0_combout ;
wire \read_data_valid~1_combout ;
wire \read_data_valid~2_combout ;
wire \read_data_valid~3_combout ;
wire \read_data_valid~q ;
wire \Equal3~5_combout ;
wire \dr_data_out[2]~14_combout ;
wire \dr_data_out[2]~15_combout ;
wire \dr_data_out~16_combout ;
wire \dr_data_out[2]~9_combout ;
wire \dr_data_out[2]~19_combout ;
wire \dr_data_out~39_combout ;
wire \dr_data_out[7]~10_combout ;
wire \dr_data_out[7]~36_combout ;
wire \dr_data_out[7]~40_combout ;
wire \dr_data_out[7]~37_combout ;
wire \dr_data_out[0]~38_combout ;
wire \dr_data_out[7]~q ;
wire \dr_data_out~34_combout ;
wire \dr_data_out~24_combout ;
wire \dr_data_out~35_combout ;
wire \dr_data_out[6]~q ;
wire \dr_data_out[5]~28_combout ;
wire \dr_data_out[5]~29_combout ;
wire \dr_data_out[5]~30_combout ;
wire \dr_data_out[5]~31_combout ;
wire \dr_data_out[5]~32_combout ;
wire \dr_data_out[5]~33_combout ;
wire \dr_data_out[5]~q ;
wire \dr_data_out~26_combout ;
wire \dr_data_out~27_combout ;
wire \dr_data_out[4]~q ;
wire \dr_data_out~23_combout ;
wire \dr_data_out~25_combout ;
wire \dr_data_out[3]~q ;
wire \dr_data_out~21_combout ;
wire \dr_data_out~22_combout ;
wire \dr_data_out[2]~q ;
wire \dr_data_out~17_combout ;
wire \dr_data_out~20_combout ;
wire \dr_data_out[1]~q ;
wire \dr_data_out~8_combout ;
wire \Selector41~2_combout ;
wire \Selector41~3_combout ;
wire \Selector41~4_combout ;
wire \dr_data_out[0]~0_combout ;
wire \dr_data_out[0]~q ;
wire \Mux0~0_combout ;
wire \Equal14~1_combout ;
wire \dr_info[8]~11_combout ;
wire \dr_info[8]~q ;
wire \dr_info~10_combout ;
wire \dr_info[0]~12_combout ;
wire \dr_info[7]~q ;
wire \dr_info~9_combout ;
wire \dr_info[6]~q ;
wire \dr_info~8_combout ;
wire \dr_info[5]~q ;
wire \dr_info~7_combout ;
wire \dr_info[4]~q ;
wire \dr_info~6_combout ;
wire \dr_info[3]~q ;
wire \dr_info~5_combout ;
wire \dr_info[2]~q ;
wire \dr_info~4_combout ;
wire \dr_info[1]~q ;
wire \dr_info~3_combout ;
wire \dr_info[0]~q ;
wire \Mux0~1_combout ;
wire \idle_inserter_source_ready~2_combout ;
wire \idle_inserter_source_ready~3_combout ;
wire \idle_inserter_source_ready~4_combout ;
wire \idle_inserter_source_ready~5_combout ;
wire \idle_inserter_source_ready~6_combout ;
wire \idle_inserter_source_ready~7_combout ;
wire \dr_data_in[1]~0_combout ;
wire \dr_data_in[7]~q ;
wire \dr_data_in[6]~q ;
wire \dr_data_in[5]~q ;
wire \dr_data_in[4]~q ;
wire \Add4~0_combout ;
wire \valid_write_data_length_byte_counter~0_combout ;
wire \decode_header_2~0_combout ;
wire \decode_header_2~1_combout ;
wire \decode_header_2~2_combout ;
wire \decode_header_2~q ;
wire \valid_write_data_length_byte_counter[5]~1_combout ;
wire \valid_write_data_length_byte_counter[0]~2_combout ;
wire \valid_write_data_length_byte_counter[0]~q ;
wire \Add4~1 ;
wire \Add4~2_combout ;
wire \valid_write_data_length_byte_counter~3_combout ;
wire \valid_write_data_length_byte_counter[1]~q ;
wire \Add4~3 ;
wire \Add4~4_combout ;
wire \valid_write_data_length_byte_counter~4_combout ;
wire \valid_write_data_length_byte_counter[2]~q ;
wire \Add4~5 ;
wire \Add4~6_combout ;
wire \valid_write_data_length_byte_counter~5_combout ;
wire \valid_write_data_length_byte_counter[3]~q ;
wire \Equal13~0_combout ;
wire \Add4~7 ;
wire \Add4~8_combout ;
wire \valid_write_data_length_byte_counter~6_combout ;
wire \valid_write_data_length_byte_counter[4]~q ;
wire \Add4~9 ;
wire \Add4~10_combout ;
wire \valid_write_data_length_byte_counter~7_combout ;
wire \valid_write_data_length_byte_counter[5]~q ;
wire \Add4~11 ;
wire \Add4~12_combout ;
wire \valid_write_data_length_byte_counter~8_combout ;
wire \valid_write_data_length_byte_counter[6]~q ;
wire \Add4~13 ;
wire \Add4~14_combout ;
wire \valid_write_data_length_byte_counter~9_combout ;
wire \valid_write_data_length_byte_counter[7]~q ;
wire \Equal13~1_combout ;
wire \write_data_length[0]~1_combout ;
wire \write_data_length[0]~q ;
wire \valid_write_data_length_byte_counter~10_combout ;
wire \write_data_length[1]~q ;
wire \write_data_length[2]~q ;
wire \valid_write_data_length_byte_counter~11_combout ;
wire \Add4~15 ;
wire \Add4~16_combout ;
wire \valid_write_data_length_byte_counter~12_combout ;
wire \valid_write_data_length_byte_counter[8]~q ;
wire \valid_write_data_length_byte_counter~13_combout ;
wire \Add2~0_combout ;
wire \valid_write_data_length_byte_counter~14_combout ;
wire \Add4~17 ;
wire \Add4~18_combout ;
wire \valid_write_data_length_byte_counter~15_combout ;
wire \valid_write_data_length_byte_counter[9]~q ;
wire \Add2~1 ;
wire \Add2~2_combout ;
wire \valid_write_data_length_byte_counter~16_combout ;
wire \Add4~19 ;
wire \Add4~20_combout ;
wire \valid_write_data_length_byte_counter~17_combout ;
wire \valid_write_data_length_byte_counter[10]~q ;
wire \Add4~21 ;
wire \Add4~22_combout ;
wire \Add2~3 ;
wire \Add2~4_combout ;
wire \valid_write_data_length_byte_counter~18_combout ;
wire \valid_write_data_length_byte_counter~19_combout ;
wire \valid_write_data_length_byte_counter[11]~q ;
wire \Equal13~2_combout ;
wire \Add2~5 ;
wire \Add2~6_combout ;
wire \valid_write_data_length_byte_counter~20_combout ;
wire \Add4~23 ;
wire \Add4~24_combout ;
wire \valid_write_data_length_byte_counter~21_combout ;
wire \valid_write_data_length_byte_counter[12]~q ;
wire \Add2~7 ;
wire \Add2~8_combout ;
wire \valid_write_data_length_byte_counter~22_combout ;
wire \Add4~25 ;
wire \Add4~26_combout ;
wire \valid_write_data_length_byte_counter~23_combout ;
wire \valid_write_data_length_byte_counter[13]~q ;
wire \Add2~9 ;
wire \Add2~10_combout ;
wire \valid_write_data_length_byte_counter~24_combout ;
wire \valid_write_data_length_byte_counter~25_combout ;
wire \Add4~27 ;
wire \Add4~28_combout ;
wire \valid_write_data_length_byte_counter~26_combout ;
wire \valid_write_data_length_byte_counter[14]~q ;
wire \Add4~29 ;
wire \Add4~30_combout ;
wire \Add2~11 ;
wire \Add2~12_combout ;
wire \valid_write_data_length_byte_counter~27_combout ;
wire \valid_write_data_length_byte_counter~28_combout ;
wire \valid_write_data_length_byte_counter[15]~q ;
wire \Equal13~3_combout ;
wire \Equal13~4_combout ;
wire \Add4~31 ;
wire \Add4~32_combout ;
wire \Add2~13 ;
wire \Add2~14_combout ;
wire \valid_write_data_length_byte_counter~29_combout ;
wire \valid_write_data_length_byte_counter~30_combout ;
wire \valid_write_data_length_byte_counter[16]~q ;
wire \Add4~33 ;
wire \Add4~34_combout ;
wire \Add2~15 ;
wire \Add2~16_combout ;
wire \valid_write_data_length_byte_counter~31_combout ;
wire \valid_write_data_length_byte_counter~32_combout ;
wire \valid_write_data_length_byte_counter[17]~q ;
wire \Add2~17 ;
wire \Add2~18_combout ;
wire \valid_write_data_length_byte_counter~33_combout ;
wire \Add4~35 ;
wire \Add4~36_combout ;
wire \valid_write_data_length_byte_counter~34_combout ;
wire \valid_write_data_length_byte_counter[18]~q ;
wire \Equal13~5_combout ;
wire \write_data_valid~q ;
wire \write_data_bit_counter~0_combout ;
wire \write_data_bit_counter[0]~1_combout ;
wire \write_data_bit_counter[0]~q ;
wire \write_data_bit_counter~2_combout ;
wire \write_data_bit_counter[1]~q ;
wire \Add3~0_combout ;
wire \write_data_bit_counter~3_combout ;
wire \write_data_bit_counter[2]~q ;
wire \always2~0_combout ;
wire \idle_remover_sink_data[0]~0_combout ;
wire \dr_data_in[3]~q ;
wire \dr_data_in[2]~q ;
wire \dr_data_in[1]~q ;


ADC_altera_avalon_st_idle_inserter idle_inserter(
	.data1_0(data1_0),
	.data1_2(data1_2),
	.data1_1(data1_1),
	.data1_6(data1_6),
	.data1_7(data1_7),
	.data1_5(data1_5),
	.data1_3(data1_3),
	.data1_4(data1_4),
	.out_data(out_data),
	.out_data1(\idle_inserter|out_data~3_combout ),
	.full1(full1),
	.reset_n(reset_n),
	.idle_inserter_source_ready(idle_inserter_source_ready1),
	.in_ready(sink_ready),
	.out_data2(\idle_inserter|out_data~4_combout ),
	.clk(altera_internal_jtag));

ADC_altera_avalon_st_idle_remover idle_remover(
	.reset_n(reset_n),
	.idle_remover_sink_data_3(idle_remover_sink_data_3),
	.idle_remover_sink_valid(\idle_remover_sink_valid~q ),
	.idle_remover_sink_data_7(idle_remover_sink_data_7),
	.idle_remover_sink_data_6(idle_remover_sink_data_6),
	.idle_remover_sink_data_4(idle_remover_sink_data_4),
	.idle_remover_sink_data_5(\idle_remover_sink_data[5]~q ),
	.idle_remover_sink_data_1(idle_remover_sink_data_1),
	.idle_remover_sink_data_0(idle_remover_sink_data_0),
	.idle_remover_sink_data_2(idle_remover_sink_data_2),
	.out_data_5(out_data_5),
	.out_valid1(out_valid),
	.clk(altera_internal_jtag));

ADC_altera_std_synchronizer_3 clock_sense_reset_n_synchronizer(
	.dreg_6(\clock_sense_reset_n_synchronizer|dreg[6]~q ),
	.reset_n(\clock_sense_reset_n~q ),
	.clk(clk_clk));

ADC_altera_std_synchronizer_5 clock_to_sample_div2_synchronizer(
	.dreg_1(\clock_to_sample_div2_synchronizer|dreg[1]~q ),
	.din(\clock_to_sample_div2~q ),
	.clk(altera_internal_jtag));

ADC_altera_std_synchronizer_6 reset_to_sample_synchronizer(
	.dreg_1(\reset_to_sample_synchronizer|dreg[1]~q ),
	.din(altera_reset_synchronizer_int_chain_out),
	.clk(altera_internal_jtag));

ADC_altera_std_synchronizer_4 clock_sensor_synchronizer(
	.dreg_1(\clock_sensor_synchronizer|dreg[1]~q ),
	.din(\clock_sensor~q ),
	.clk(altera_internal_jtag));

dffeas clock_to_sample_div2(
	.clk(clk_clk),
	.d(\clock_to_sample_div2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\clock_to_sample_div2~q ),
	.prn(vcc));
defparam clock_to_sample_div2.is_wysiwyg = "true";
defparam clock_to_sample_div2.power_up = "low";

dffeas clock_sensor(
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(\clock_sense_reset_n_synchronizer|dreg[6]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\clock_sensor~q ),
	.prn(vcc));
defparam clock_sensor.is_wysiwyg = "true";
defparam clock_sensor.power_up = "low";

dffeas clock_sense_reset_n(
	.clk(altera_internal_jtag),
	.d(virtual_state_udr),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal14~2_combout ),
	.q(\clock_sense_reset_n~q ),
	.prn(vcc));
defparam clock_sense_reset_n.is_wysiwyg = "true";
defparam clock_sense_reset_n.power_up = "low";

dffeas idle_remover_sink_valid(
	.clk(altera_internal_jtag),
	.d(\idle_remover_sink_data[0]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\idle_remover_sink_valid~q ),
	.prn(vcc));
defparam idle_remover_sink_valid.is_wysiwyg = "true";
defparam idle_remover_sink_valid.power_up = "low";

dffeas \idle_remover_sink_data[5] (
	.clk(altera_internal_jtag),
	.d(\dr_data_in[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idle_remover_sink_data[0]~0_combout ),
	.q(\idle_remover_sink_data[5]~q ),
	.prn(vcc));
defparam \idle_remover_sink_data[5] .is_wysiwyg = "true";
defparam \idle_remover_sink_data[5] .power_up = "low";

fiftyfivenm_lcell_comb \clock_to_sample_div2~0 (
	.dataa(\clock_to_sample_div2~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\clock_to_sample_div2~0_combout ),
	.cout());
defparam \clock_to_sample_div2~0 .lut_mask = 16'h5555;
defparam \clock_to_sample_div2~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \tdo~1 (
	.dataa(virtual_state_sdr),
	.datab(\tdo~0_combout ),
	.datac(\Mux0~1_combout ),
	.datad(irf_reg_2_1),
	.cin(gnd),
	.combout(tdo),
	.cout());
defparam \tdo~1 .lut_mask = 16'hFDFF;
defparam \tdo~1 .sum_lutc_input = "datac";

dffeas idle_inserter_source_ready(
	.clk(altera_internal_jtag),
	.d(\idle_inserter_source_ready~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(idle_inserter_source_ready1),
	.prn(vcc));
defparam idle_inserter_source_ready.is_wysiwyg = "true";
defparam idle_inserter_source_ready.power_up = "low";

dffeas \idle_remover_sink_data[3] (
	.clk(altera_internal_jtag),
	.d(\dr_data_in[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idle_remover_sink_data[0]~0_combout ),
	.q(idle_remover_sink_data_3),
	.prn(vcc));
defparam \idle_remover_sink_data[3] .is_wysiwyg = "true";
defparam \idle_remover_sink_data[3] .power_up = "low";

dffeas \idle_remover_sink_data[7] (
	.clk(altera_internal_jtag),
	.d(altera_internal_jtag1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idle_remover_sink_data[0]~0_combout ),
	.q(idle_remover_sink_data_7),
	.prn(vcc));
defparam \idle_remover_sink_data[7] .is_wysiwyg = "true";
defparam \idle_remover_sink_data[7] .power_up = "low";

dffeas \idle_remover_sink_data[6] (
	.clk(altera_internal_jtag),
	.d(\dr_data_in[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idle_remover_sink_data[0]~0_combout ),
	.q(idle_remover_sink_data_6),
	.prn(vcc));
defparam \idle_remover_sink_data[6] .is_wysiwyg = "true";
defparam \idle_remover_sink_data[6] .power_up = "low";

dffeas \idle_remover_sink_data[4] (
	.clk(altera_internal_jtag),
	.d(\dr_data_in[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idle_remover_sink_data[0]~0_combout ),
	.q(idle_remover_sink_data_4),
	.prn(vcc));
defparam \idle_remover_sink_data[4] .is_wysiwyg = "true";
defparam \idle_remover_sink_data[4] .power_up = "low";

dffeas \idle_remover_sink_data[1] (
	.clk(altera_internal_jtag),
	.d(\dr_data_in[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idle_remover_sink_data[0]~0_combout ),
	.q(idle_remover_sink_data_1),
	.prn(vcc));
defparam \idle_remover_sink_data[1] .is_wysiwyg = "true";
defparam \idle_remover_sink_data[1] .power_up = "low";

dffeas \idle_remover_sink_data[0] (
	.clk(altera_internal_jtag),
	.d(\dr_data_in[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idle_remover_sink_data[0]~0_combout ),
	.q(idle_remover_sink_data_0),
	.prn(vcc));
defparam \idle_remover_sink_data[0] .is_wysiwyg = "true";
defparam \idle_remover_sink_data[0] .power_up = "low";

dffeas \idle_remover_sink_data[2] (
	.clk(altera_internal_jtag),
	.d(\dr_data_in[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\idle_remover_sink_data[0]~0_combout ),
	.q(idle_remover_sink_data_2),
	.prn(vcc));
defparam \idle_remover_sink_data[2] .is_wysiwyg = "true";
defparam \idle_remover_sink_data[2] .power_up = "low";

fiftyfivenm_lcell_comb \dr_loopback~0 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(state_4),
	.datac(altera_internal_jtag1),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\dr_loopback~0_combout ),
	.cout());
defparam \dr_loopback~0 .lut_mask = 16'hFEFF;
defparam \dr_loopback~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dr_info[4]~2 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(state_4),
	.datac(state_3),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\dr_info[4]~2_combout ),
	.cout());
defparam \dr_info[4]~2 .lut_mask = 16'hFEFF;
defparam \dr_info[4]~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dr_control[0]~1 (
	.dataa(irf_reg_2_1),
	.datab(\dr_info[4]~2_combout ),
	.datac(irf_reg_0_1),
	.datad(irf_reg_1_1),
	.cin(gnd),
	.combout(\dr_control[0]~1_combout ),
	.cout());
defparam \dr_control[0]~1 .lut_mask = 16'hEFFF;
defparam \dr_control[0]~1 .sum_lutc_input = "datac";

dffeas \dr_control[8] (
	.clk(altera_internal_jtag),
	.d(\dr_loopback~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dr_control[0]~1_combout ),
	.q(\dr_control[8]~q ),
	.prn(vcc));
defparam \dr_control[8] .is_wysiwyg = "true";
defparam \dr_control[8] .power_up = "low";

fiftyfivenm_lcell_comb \dr_control~8 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(state_4),
	.datac(\dr_control[8]~q ),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\dr_control~8_combout ),
	.cout());
defparam \dr_control~8 .lut_mask = 16'hFEFF;
defparam \dr_control~8 .sum_lutc_input = "datac";

dffeas \dr_control[7] (
	.clk(altera_internal_jtag),
	.d(\dr_control~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dr_control[0]~1_combout ),
	.q(\dr_control[7]~q ),
	.prn(vcc));
defparam \dr_control[7] .is_wysiwyg = "true";
defparam \dr_control[7] .power_up = "low";

fiftyfivenm_lcell_comb \dr_control~7 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(state_4),
	.datac(\dr_control[7]~q ),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\dr_control~7_combout ),
	.cout());
defparam \dr_control~7 .lut_mask = 16'hFEFF;
defparam \dr_control~7 .sum_lutc_input = "datac";

dffeas \dr_control[6] (
	.clk(altera_internal_jtag),
	.d(\dr_control~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dr_control[0]~1_combout ),
	.q(\dr_control[6]~q ),
	.prn(vcc));
defparam \dr_control[6] .is_wysiwyg = "true";
defparam \dr_control[6] .power_up = "low";

fiftyfivenm_lcell_comb \dr_control~6 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(state_4),
	.datac(\dr_control[6]~q ),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\dr_control~6_combout ),
	.cout());
defparam \dr_control~6 .lut_mask = 16'hFEFF;
defparam \dr_control~6 .sum_lutc_input = "datac";

dffeas \dr_control[5] (
	.clk(altera_internal_jtag),
	.d(\dr_control~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dr_control[0]~1_combout ),
	.q(\dr_control[5]~q ),
	.prn(vcc));
defparam \dr_control[5] .is_wysiwyg = "true";
defparam \dr_control[5] .power_up = "low";

fiftyfivenm_lcell_comb \dr_control~5 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(state_4),
	.datac(\dr_control[5]~q ),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\dr_control~5_combout ),
	.cout());
defparam \dr_control~5 .lut_mask = 16'hFEFF;
defparam \dr_control~5 .sum_lutc_input = "datac";

dffeas \dr_control[4] (
	.clk(altera_internal_jtag),
	.d(\dr_control~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dr_control[0]~1_combout ),
	.q(\dr_control[4]~q ),
	.prn(vcc));
defparam \dr_control[4] .is_wysiwyg = "true";
defparam \dr_control[4] .power_up = "low";

fiftyfivenm_lcell_comb \dr_control~4 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(state_4),
	.datac(\dr_control[4]~q ),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\dr_control~4_combout ),
	.cout());
defparam \dr_control~4 .lut_mask = 16'hFEFF;
defparam \dr_control~4 .sum_lutc_input = "datac";

dffeas \dr_control[3] (
	.clk(altera_internal_jtag),
	.d(\dr_control~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dr_control[0]~1_combout ),
	.q(\dr_control[3]~q ),
	.prn(vcc));
defparam \dr_control[3] .is_wysiwyg = "true";
defparam \dr_control[3] .power_up = "low";

fiftyfivenm_lcell_comb \dr_control~3 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(state_4),
	.datac(\dr_control[3]~q ),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\dr_control~3_combout ),
	.cout());
defparam \dr_control~3 .lut_mask = 16'hFEFF;
defparam \dr_control~3 .sum_lutc_input = "datac";

dffeas \dr_control[2] (
	.clk(altera_internal_jtag),
	.d(\dr_control~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dr_control[0]~1_combout ),
	.q(\dr_control[2]~q ),
	.prn(vcc));
defparam \dr_control[2] .is_wysiwyg = "true";
defparam \dr_control[2] .power_up = "low";

fiftyfivenm_lcell_comb \dr_control~2 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(state_4),
	.datac(\dr_control[2]~q ),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\dr_control~2_combout ),
	.cout());
defparam \dr_control~2 .lut_mask = 16'hFEFF;
defparam \dr_control~2 .sum_lutc_input = "datac";

dffeas \dr_control[1] (
	.clk(altera_internal_jtag),
	.d(\dr_control~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dr_control[0]~1_combout ),
	.q(\dr_control[1]~q ),
	.prn(vcc));
defparam \dr_control[1] .is_wysiwyg = "true";
defparam \dr_control[1] .power_up = "low";

fiftyfivenm_lcell_comb \dr_control~0 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(state_4),
	.datac(\dr_control[1]~q ),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\dr_control~0_combout ),
	.cout());
defparam \dr_control~0 .lut_mask = 16'hFEFF;
defparam \dr_control~0 .sum_lutc_input = "datac";

dffeas \dr_control[0] (
	.clk(altera_internal_jtag),
	.d(\dr_control~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dr_control[0]~1_combout ),
	.q(\dr_control[0]~q ),
	.prn(vcc));
defparam \dr_control[0] .is_wysiwyg = "true";
defparam \dr_control[0] .power_up = "low";

fiftyfivenm_lcell_comb \tdo~0 (
	.dataa(\dr_control[0]~q ),
	.datab(irf_reg_2_1),
	.datac(irf_reg_0_1),
	.datad(irf_reg_1_1),
	.cin(gnd),
	.combout(\tdo~0_combout ),
	.cout());
defparam \tdo~0 .lut_mask = 16'hEFFF;
defparam \tdo~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dr_debug~3 (
	.dataa(\dr_debug[2]~q ),
	.datab(\clock_sensor_synchronizer|dreg[1]~q ),
	.datac(virtual_state_cdr),
	.datad(virtual_state_sdr),
	.cin(gnd),
	.combout(\dr_debug~3_combout ),
	.cout());
defparam \dr_debug~3 .lut_mask = 16'hFFAC;
defparam \dr_debug~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Equal14~2 (
	.dataa(irf_reg_1_1),
	.datab(gnd),
	.datac(irf_reg_2_1),
	.datad(irf_reg_0_1),
	.cin(gnd),
	.combout(\Equal14~2_combout ),
	.cout());
defparam \Equal14~2 .lut_mask = 16'hAFFF;
defparam \Equal14~2 .sum_lutc_input = "datac";

dffeas \dr_debug[2] (
	.clk(altera_internal_jtag),
	.d(\dr_debug~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal14~2_combout ),
	.q(\dr_debug[2]~q ),
	.prn(vcc));
defparam \dr_debug[2] .is_wysiwyg = "true";
defparam \dr_debug[2] .power_up = "low";

fiftyfivenm_lcell_comb \dr_debug~2 (
	.dataa(\dr_debug[2]~q ),
	.datab(\clock_to_sample_div2_synchronizer|dreg[1]~q ),
	.datac(gnd),
	.datad(virtual_state_sdr),
	.cin(gnd),
	.combout(\dr_debug~2_combout ),
	.cout());
defparam \dr_debug~2 .lut_mask = 16'hAACC;
defparam \dr_debug~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dr_debug[0]~1 (
	.dataa(irf_reg_1_1),
	.datab(\dr_info[4]~2_combout ),
	.datac(irf_reg_2_1),
	.datad(irf_reg_0_1),
	.cin(gnd),
	.combout(\dr_debug[0]~1_combout ),
	.cout());
defparam \dr_debug[0]~1 .lut_mask = 16'hEFFF;
defparam \dr_debug[0]~1 .sum_lutc_input = "datac";

dffeas \dr_debug[1] (
	.clk(altera_internal_jtag),
	.d(\dr_debug~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dr_debug[0]~1_combout ),
	.q(\dr_debug[1]~q ),
	.prn(vcc));
defparam \dr_debug[1] .is_wysiwyg = "true";
defparam \dr_debug[1] .power_up = "low";

fiftyfivenm_lcell_comb \dr_debug~0 (
	.dataa(\dr_debug[1]~q ),
	.datab(\reset_to_sample_synchronizer|dreg[1]~q ),
	.datac(gnd),
	.datad(virtual_state_sdr),
	.cin(gnd),
	.combout(\dr_debug~0_combout ),
	.cout());
defparam \dr_debug~0 .lut_mask = 16'hAACC;
defparam \dr_debug~0 .sum_lutc_input = "datac";

dffeas \dr_debug[0] (
	.clk(altera_internal_jtag),
	.d(\dr_debug~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dr_debug[0]~1_combout ),
	.q(\dr_debug[0]~q ),
	.prn(vcc));
defparam \dr_debug[0] .is_wysiwyg = "true";
defparam \dr_debug[0] .power_up = "low";

fiftyfivenm_lcell_comb \dr_loopback~1 (
	.dataa(irf_reg_0_1),
	.datab(gnd),
	.datac(irf_reg_2_1),
	.datad(irf_reg_1_1),
	.cin(gnd),
	.combout(\dr_loopback~1_combout ),
	.cout());
defparam \dr_loopback~1 .lut_mask = 16'hAFFF;
defparam \dr_loopback~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dr_loopback~2 (
	.dataa(\dr_loopback~0_combout ),
	.datab(\dr_loopback~q ),
	.datac(\dr_info[4]~2_combout ),
	.datad(\dr_loopback~1_combout ),
	.cin(gnd),
	.combout(\dr_loopback~2_combout ),
	.cout());
defparam \dr_loopback~2 .lut_mask = 16'hEFFE;
defparam \dr_loopback~2 .sum_lutc_input = "datac";

dffeas dr_loopback(
	.clk(altera_internal_jtag),
	.d(\dr_loopback~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dr_loopback~q ),
	.prn(vcc));
defparam dr_loopback.is_wysiwyg = "true";
defparam dr_loopback.power_up = "low";

fiftyfivenm_lcell_comb \read_data_all_valid~0 (
	.dataa(\read_data_all_valid~q ),
	.datab(virtual_ir_scan_reg),
	.datac(splitter_nodes_receive_0_3),
	.datad(state_3),
	.cin(gnd),
	.combout(\read_data_all_valid~0_combout ),
	.cout());
defparam \read_data_all_valid~0 .lut_mask = 16'hEFFF;
defparam \read_data_all_valid~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Equal14~0 (
	.dataa(gnd),
	.datab(irf_reg_2_1),
	.datac(irf_reg_0_1),
	.datad(irf_reg_1_1),
	.cin(gnd),
	.combout(\Equal14~0_combout ),
	.cout());
defparam \Equal14~0 .lut_mask = 16'h3FFF;
defparam \Equal14~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \offset[7]~0 (
	.dataa(irf_reg_2_1),
	.datab(virtual_state_udr),
	.datac(irf_reg_0_1),
	.datad(irf_reg_1_1),
	.cin(gnd),
	.combout(\offset[7]~0_combout ),
	.cout());
defparam \offset[7]~0 .lut_mask = 16'hEFFF;
defparam \offset[7]~0 .sum_lutc_input = "datac";

dffeas \offset[2] (
	.clk(altera_internal_jtag),
	.d(\dr_control[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\offset[7]~0_combout ),
	.q(\offset[2]~q ),
	.prn(vcc));
defparam \offset[2] .is_wysiwyg = "true";
defparam \offset[2] .power_up = "low";

dffeas \offset[1] (
	.clk(altera_internal_jtag),
	.d(\dr_control[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\offset[7]~0_combout ),
	.q(\offset[1]~q ),
	.prn(vcc));
defparam \offset[1] .is_wysiwyg = "true";
defparam \offset[1] .power_up = "low";

dffeas \offset[0] (
	.clk(altera_internal_jtag),
	.d(\dr_control[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\offset[7]~0_combout ),
	.q(\offset[0]~q ),
	.prn(vcc));
defparam \offset[0] .is_wysiwyg = "true";
defparam \offset[0] .power_up = "low";

fiftyfivenm_lcell_comb \Equal6~0 (
	.dataa(gnd),
	.datab(\offset[2]~q ),
	.datac(\offset[1]~q ),
	.datad(\offset[0]~q ),
	.cin(gnd),
	.combout(\Equal6~0_combout ),
	.cout());
defparam \Equal6~0 .lut_mask = 16'h3FFF;
defparam \Equal6~0 .sum_lutc_input = "datac";

dffeas \offset[3] (
	.clk(altera_internal_jtag),
	.d(\dr_control[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\offset[7]~0_combout ),
	.q(\offset[3]~q ),
	.prn(vcc));
defparam \offset[3] .is_wysiwyg = "true";
defparam \offset[3] .power_up = "low";

dffeas \offset[4] (
	.clk(altera_internal_jtag),
	.d(\dr_control[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\offset[7]~0_combout ),
	.q(\offset[4]~q ),
	.prn(vcc));
defparam \offset[4] .is_wysiwyg = "true";
defparam \offset[4] .power_up = "low";

dffeas \offset[5] (
	.clk(altera_internal_jtag),
	.d(\dr_control[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\offset[7]~0_combout ),
	.q(\offset[5]~q ),
	.prn(vcc));
defparam \offset[5] .is_wysiwyg = "true";
defparam \offset[5] .power_up = "low";

dffeas \offset[6] (
	.clk(altera_internal_jtag),
	.d(\dr_control[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\offset[7]~0_combout ),
	.q(\offset[6]~q ),
	.prn(vcc));
defparam \offset[6] .is_wysiwyg = "true";
defparam \offset[6] .power_up = "low";

fiftyfivenm_lcell_comb \Equal6~1 (
	.dataa(\offset[3]~q ),
	.datab(\offset[4]~q ),
	.datac(\offset[5]~q ),
	.datad(\offset[6]~q ),
	.cin(gnd),
	.combout(\Equal6~1_combout ),
	.cout());
defparam \Equal6~1 .lut_mask = 16'h7FFF;
defparam \Equal6~1 .sum_lutc_input = "datac";

dffeas \offset[7] (
	.clk(altera_internal_jtag),
	.d(\dr_control[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\offset[7]~0_combout ),
	.q(\offset[7]~q ),
	.prn(vcc));
defparam \offset[7] .is_wysiwyg = "true";
defparam \offset[7] .power_up = "low";

fiftyfivenm_lcell_comb \Equal6~2 (
	.dataa(\Equal6~0_combout ),
	.datab(\Equal6~1_combout ),
	.datac(gnd),
	.datad(\offset[7]~q ),
	.cin(gnd),
	.combout(\Equal6~2_combout ),
	.cout());
defparam \Equal6~2 .lut_mask = 16'hEEFF;
defparam \Equal6~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \write_state~22 (
	.dataa(\Equal6~0_combout ),
	.datab(\Equal6~1_combout ),
	.datac(\offset[7]~q ),
	.datad(\write_state~17_combout ),
	.cin(gnd),
	.combout(\write_state~22_combout ),
	.cout());
defparam \write_state~22 .lut_mask = 16'hEFFF;
defparam \write_state~22 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \write_state~19 (
	.dataa(virtual_state_cdr),
	.datab(\write_state~17_combout ),
	.datac(gnd),
	.datad(\Equal14~0_combout ),
	.cin(gnd),
	.combout(\write_state~19_combout ),
	.cout());
defparam \write_state~19 .lut_mask = 16'hFF77;
defparam \write_state~19 .sum_lutc_input = "datac";

dffeas \write_state.ST_BYPASS (
	.clk(altera_internal_jtag),
	.d(\write_state~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_state~19_combout ),
	.q(\write_state.ST_BYPASS~q ),
	.prn(vcc));
defparam \write_state.ST_BYPASS .is_wysiwyg = "true";
defparam \write_state.ST_BYPASS .power_up = "low";

fiftyfivenm_lcell_comb \bypass_bit_counter[0]~8 (
	.dataa(\bypass_bit_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\bypass_bit_counter[0]~8_combout ),
	.cout(\bypass_bit_counter[0]~9 ));
defparam \bypass_bit_counter[0]~8 .lut_mask = 16'h55AA;
defparam \bypass_bit_counter[0]~8 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \bypass_bit_counter~12 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(state_4),
	.datac(virtual_ir_scan_reg),
	.datad(\write_state.ST_BYPASS~q ),
	.cin(gnd),
	.combout(\bypass_bit_counter~12_combout ),
	.cout());
defparam \bypass_bit_counter~12 .lut_mask = 16'hFFF7;
defparam \bypass_bit_counter~12 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \bypass_bit_counter[0]~13 (
	.dataa(\Equal14~0_combout ),
	.datab(virtual_state_sdr),
	.datac(\write_state.ST_BYPASS~q ),
	.datad(virtual_state_cdr),
	.cin(gnd),
	.combout(\bypass_bit_counter[0]~13_combout ),
	.cout());
defparam \bypass_bit_counter[0]~13 .lut_mask = 16'hBFFF;
defparam \bypass_bit_counter[0]~13 .sum_lutc_input = "datac";

dffeas \bypass_bit_counter[0] (
	.clk(altera_internal_jtag),
	.d(\bypass_bit_counter[0]~8_combout ),
	.asdata(\offset[0]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\bypass_bit_counter~12_combout ),
	.ena(\bypass_bit_counter[0]~13_combout ),
	.q(\bypass_bit_counter[0]~q ),
	.prn(vcc));
defparam \bypass_bit_counter[0] .is_wysiwyg = "true";
defparam \bypass_bit_counter[0] .power_up = "low";

fiftyfivenm_lcell_comb \bypass_bit_counter[1]~10 (
	.dataa(\bypass_bit_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\bypass_bit_counter[0]~9 ),
	.combout(\bypass_bit_counter[1]~10_combout ),
	.cout(\bypass_bit_counter[1]~11 ));
defparam \bypass_bit_counter[1]~10 .lut_mask = 16'h5A5F;
defparam \bypass_bit_counter[1]~10 .sum_lutc_input = "cin";

dffeas \bypass_bit_counter[1] (
	.clk(altera_internal_jtag),
	.d(\bypass_bit_counter[1]~10_combout ),
	.asdata(\offset[1]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\bypass_bit_counter~12_combout ),
	.ena(\bypass_bit_counter[0]~13_combout ),
	.q(\bypass_bit_counter[1]~q ),
	.prn(vcc));
defparam \bypass_bit_counter[1] .is_wysiwyg = "true";
defparam \bypass_bit_counter[1] .power_up = "low";

fiftyfivenm_lcell_comb \bypass_bit_counter[2]~14 (
	.dataa(\bypass_bit_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\bypass_bit_counter[1]~11 ),
	.combout(\bypass_bit_counter[2]~14_combout ),
	.cout(\bypass_bit_counter[2]~15 ));
defparam \bypass_bit_counter[2]~14 .lut_mask = 16'h5AAF;
defparam \bypass_bit_counter[2]~14 .sum_lutc_input = "cin";

dffeas \bypass_bit_counter[2] (
	.clk(altera_internal_jtag),
	.d(\bypass_bit_counter[2]~14_combout ),
	.asdata(\offset[2]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\bypass_bit_counter~12_combout ),
	.ena(\bypass_bit_counter[0]~13_combout ),
	.q(\bypass_bit_counter[2]~q ),
	.prn(vcc));
defparam \bypass_bit_counter[2] .is_wysiwyg = "true";
defparam \bypass_bit_counter[2] .power_up = "low";

fiftyfivenm_lcell_comb \write_state~14 (
	.dataa(\write_state.ST_BYPASS~q ),
	.datab(\bypass_bit_counter[1]~q ),
	.datac(\bypass_bit_counter[2]~q ),
	.datad(\bypass_bit_counter[0]~q ),
	.cin(gnd),
	.combout(\write_state~14_combout ),
	.cout());
defparam \write_state~14 .lut_mask = 16'hFEFF;
defparam \write_state~14 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \bypass_bit_counter[3]~16 (
	.dataa(\bypass_bit_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\bypass_bit_counter[2]~15 ),
	.combout(\bypass_bit_counter[3]~16_combout ),
	.cout(\bypass_bit_counter[3]~17 ));
defparam \bypass_bit_counter[3]~16 .lut_mask = 16'h5A5F;
defparam \bypass_bit_counter[3]~16 .sum_lutc_input = "cin";

dffeas \bypass_bit_counter[3] (
	.clk(altera_internal_jtag),
	.d(\bypass_bit_counter[3]~16_combout ),
	.asdata(\offset[3]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\bypass_bit_counter~12_combout ),
	.ena(\bypass_bit_counter[0]~13_combout ),
	.q(\bypass_bit_counter[3]~q ),
	.prn(vcc));
defparam \bypass_bit_counter[3] .is_wysiwyg = "true";
defparam \bypass_bit_counter[3] .power_up = "low";

fiftyfivenm_lcell_comb \bypass_bit_counter[4]~18 (
	.dataa(\bypass_bit_counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\bypass_bit_counter[3]~17 ),
	.combout(\bypass_bit_counter[4]~18_combout ),
	.cout(\bypass_bit_counter[4]~19 ));
defparam \bypass_bit_counter[4]~18 .lut_mask = 16'h5AAF;
defparam \bypass_bit_counter[4]~18 .sum_lutc_input = "cin";

dffeas \bypass_bit_counter[4] (
	.clk(altera_internal_jtag),
	.d(\bypass_bit_counter[4]~18_combout ),
	.asdata(\offset[4]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\bypass_bit_counter~12_combout ),
	.ena(\bypass_bit_counter[0]~13_combout ),
	.q(\bypass_bit_counter[4]~q ),
	.prn(vcc));
defparam \bypass_bit_counter[4] .is_wysiwyg = "true";
defparam \bypass_bit_counter[4] .power_up = "low";

fiftyfivenm_lcell_comb \bypass_bit_counter[5]~20 (
	.dataa(\bypass_bit_counter[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\bypass_bit_counter[4]~19 ),
	.combout(\bypass_bit_counter[5]~20_combout ),
	.cout(\bypass_bit_counter[5]~21 ));
defparam \bypass_bit_counter[5]~20 .lut_mask = 16'h5A5F;
defparam \bypass_bit_counter[5]~20 .sum_lutc_input = "cin";

dffeas \bypass_bit_counter[5] (
	.clk(altera_internal_jtag),
	.d(\bypass_bit_counter[5]~20_combout ),
	.asdata(\offset[5]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\bypass_bit_counter~12_combout ),
	.ena(\bypass_bit_counter[0]~13_combout ),
	.q(\bypass_bit_counter[5]~q ),
	.prn(vcc));
defparam \bypass_bit_counter[5] .is_wysiwyg = "true";
defparam \bypass_bit_counter[5] .power_up = "low";

fiftyfivenm_lcell_comb \bypass_bit_counter[6]~22 (
	.dataa(\bypass_bit_counter[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\bypass_bit_counter[5]~21 ),
	.combout(\bypass_bit_counter[6]~22_combout ),
	.cout(\bypass_bit_counter[6]~23 ));
defparam \bypass_bit_counter[6]~22 .lut_mask = 16'h5AAF;
defparam \bypass_bit_counter[6]~22 .sum_lutc_input = "cin";

dffeas \bypass_bit_counter[6] (
	.clk(altera_internal_jtag),
	.d(\bypass_bit_counter[6]~22_combout ),
	.asdata(\offset[6]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\bypass_bit_counter~12_combout ),
	.ena(\bypass_bit_counter[0]~13_combout ),
	.q(\bypass_bit_counter[6]~q ),
	.prn(vcc));
defparam \bypass_bit_counter[6] .is_wysiwyg = "true";
defparam \bypass_bit_counter[6] .power_up = "low";

fiftyfivenm_lcell_comb \bypass_bit_counter[7]~24 (
	.dataa(\bypass_bit_counter[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\bypass_bit_counter[6]~23 ),
	.combout(\bypass_bit_counter[7]~24_combout ),
	.cout());
defparam \bypass_bit_counter[7]~24 .lut_mask = 16'h5A5A;
defparam \bypass_bit_counter[7]~24 .sum_lutc_input = "cin";

dffeas \bypass_bit_counter[7] (
	.clk(altera_internal_jtag),
	.d(\bypass_bit_counter[7]~24_combout ),
	.asdata(\offset[7]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\bypass_bit_counter~12_combout ),
	.ena(\bypass_bit_counter[0]~13_combout ),
	.q(\bypass_bit_counter[7]~q ),
	.prn(vcc));
defparam \bypass_bit_counter[7] .is_wysiwyg = "true";
defparam \bypass_bit_counter[7] .power_up = "low";

fiftyfivenm_lcell_comb \write_state~15 (
	.dataa(\bypass_bit_counter[3]~q ),
	.datab(\bypass_bit_counter[4]~q ),
	.datac(\bypass_bit_counter[5]~q ),
	.datad(\bypass_bit_counter[6]~q ),
	.cin(gnd),
	.combout(\write_state~15_combout ),
	.cout());
defparam \write_state~15 .lut_mask = 16'hFFFE;
defparam \write_state~15 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \write_state~16 (
	.dataa(\write_state~14_combout ),
	.datab(\bypass_bit_counter[7]~q ),
	.datac(\write_state~15_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\write_state~16_combout ),
	.cout());
defparam \write_state~16 .lut_mask = 16'hFEFE;
defparam \write_state~16 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \write_state~18 (
	.dataa(\write_state.ST_HEADER_1~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\write_state~17_combout ),
	.cin(gnd),
	.combout(\write_state~18_combout ),
	.cout());
defparam \write_state~18 .lut_mask = 16'hAAFF;
defparam \write_state~18 .sum_lutc_input = "datac";

dffeas \write_state.ST_HEADER_2 (
	.clk(altera_internal_jtag),
	.d(\write_state~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_state~19_combout ),
	.q(\write_state.ST_HEADER_2~q ),
	.prn(vcc));
defparam \write_state.ST_HEADER_2 .is_wysiwyg = "true";
defparam \write_state.ST_HEADER_2 .power_up = "low";

fiftyfivenm_lcell_comb \write_state~21 (
	.dataa(\write_state.ST_HEADER_2~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\write_state~17_combout ),
	.cin(gnd),
	.combout(\write_state~21_combout ),
	.cout());
defparam \write_state~21 .lut_mask = 16'hAAFF;
defparam \write_state~21 .sum_lutc_input = "datac";

dffeas \write_state.ST_WRITE_DATA (
	.clk(altera_internal_jtag),
	.d(\write_state~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_state~19_combout ),
	.q(\write_state.ST_WRITE_DATA~q ),
	.prn(vcc));
defparam \write_state.ST_WRITE_DATA .is_wysiwyg = "true";
defparam \write_state.ST_WRITE_DATA .power_up = "low";

fiftyfivenm_lcell_comb \header_in_bit_counter~3 (
	.dataa(\write_state.ST_WRITE_DATA~q ),
	.datab(virtual_state_sdr),
	.datac(\header_in_bit_counter[0]~q ),
	.datad(\write_state.ST_BYPASS~q ),
	.cin(gnd),
	.combout(\header_in_bit_counter~3_combout ),
	.cout());
defparam \header_in_bit_counter~3 .lut_mask = 16'hEFFF;
defparam \header_in_bit_counter~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \header_in_bit_counter[0]~4 (
	.dataa(state_3),
	.datab(state_4),
	.datac(\write_state.ST_BYPASS~q ),
	.datad(\write_state.ST_WRITE_DATA~q ),
	.cin(gnd),
	.combout(\header_in_bit_counter[0]~4_combout ),
	.cout());
defparam \header_in_bit_counter[0]~4 .lut_mask = 16'hFEFF;
defparam \header_in_bit_counter[0]~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \header_in_bit_counter[0]~5 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(\Equal14~0_combout ),
	.datac(\header_in_bit_counter[0]~4_combout ),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\header_in_bit_counter[0]~5_combout ),
	.cout());
defparam \header_in_bit_counter[0]~5 .lut_mask = 16'hFEFF;
defparam \header_in_bit_counter[0]~5 .sum_lutc_input = "datac";

dffeas \header_in_bit_counter[0] (
	.clk(altera_internal_jtag),
	.d(\header_in_bit_counter~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\header_in_bit_counter[0]~5_combout ),
	.q(\header_in_bit_counter[0]~q ),
	.prn(vcc));
defparam \header_in_bit_counter[0] .is_wysiwyg = "true";
defparam \header_in_bit_counter[0] .power_up = "low";

fiftyfivenm_lcell_comb \header_in_bit_counter~2 (
	.dataa(virtual_state_sdr),
	.datab(\write_state.ST_BYPASS~q ),
	.datac(gnd),
	.datad(\write_state.ST_WRITE_DATA~q ),
	.cin(gnd),
	.combout(\header_in_bit_counter~2_combout ),
	.cout());
defparam \header_in_bit_counter~2 .lut_mask = 16'hDDFF;
defparam \header_in_bit_counter~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \header_in_bit_counter~6 (
	.dataa(\header_in_bit_counter[0]~q ),
	.datab(\header_in_bit_counter[1]~q ),
	.datac(gnd),
	.datad(\header_in_bit_counter~2_combout ),
	.cin(gnd),
	.combout(\header_in_bit_counter~6_combout ),
	.cout());
defparam \header_in_bit_counter~6 .lut_mask = 16'h66FF;
defparam \header_in_bit_counter~6 .sum_lutc_input = "datac";

dffeas \header_in_bit_counter[1] (
	.clk(altera_internal_jtag),
	.d(\header_in_bit_counter~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\header_in_bit_counter[0]~5_combout ),
	.q(\header_in_bit_counter[1]~q ),
	.prn(vcc));
defparam \header_in_bit_counter[1] .is_wysiwyg = "true";
defparam \header_in_bit_counter[1] .power_up = "low";

fiftyfivenm_lcell_comb \header_in_bit_counter~8 (
	.dataa(\header_in_bit_counter[0]~q ),
	.datab(\header_in_bit_counter[1]~q ),
	.datac(\header_in_bit_counter[2]~q ),
	.datad(\header_in_bit_counter~2_combout ),
	.cin(gnd),
	.combout(\header_in_bit_counter~8_combout ),
	.cout());
defparam \header_in_bit_counter~8 .lut_mask = 16'h96FF;
defparam \header_in_bit_counter~8 .sum_lutc_input = "datac";

dffeas \header_in_bit_counter[2] (
	.clk(altera_internal_jtag),
	.d(\header_in_bit_counter~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\header_in_bit_counter[0]~5_combout ),
	.q(\header_in_bit_counter[2]~q ),
	.prn(vcc));
defparam \header_in_bit_counter[2] .is_wysiwyg = "true";
defparam \header_in_bit_counter[2] .power_up = "low";

fiftyfivenm_lcell_comb \Add1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\header_in_bit_counter[0]~q ),
	.datad(\header_in_bit_counter[1]~q ),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout());
defparam \Add1~0 .lut_mask = 16'h0FFF;
defparam \Add1~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \header_in_bit_counter~7 (
	.dataa(\header_in_bit_counter[3]~q ),
	.datab(\header_in_bit_counter[2]~q ),
	.datac(\Add1~0_combout ),
	.datad(\header_in_bit_counter~2_combout ),
	.cin(gnd),
	.combout(\header_in_bit_counter~7_combout ),
	.cout());
defparam \header_in_bit_counter~7 .lut_mask = 16'h96FF;
defparam \header_in_bit_counter~7 .sum_lutc_input = "datac";

dffeas \header_in_bit_counter[3] (
	.clk(altera_internal_jtag),
	.d(\header_in_bit_counter~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\header_in_bit_counter[0]~5_combout ),
	.q(\header_in_bit_counter[3]~q ),
	.prn(vcc));
defparam \header_in_bit_counter[3] .is_wysiwyg = "true";
defparam \header_in_bit_counter[3] .power_up = "low";

fiftyfivenm_lcell_comb \read_data_length[0]~0 (
	.dataa(\header_in_bit_counter[0]~q ),
	.datab(\header_in_bit_counter[1]~q ),
	.datac(\header_in_bit_counter[2]~q ),
	.datad(\header_in_bit_counter[3]~q ),
	.cin(gnd),
	.combout(\read_data_length[0]~0_combout ),
	.cout());
defparam \read_data_length[0]~0 .lut_mask = 16'hEFFF;
defparam \read_data_length[0]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \read_data_length[0]~2 (
	.dataa(\write_state.ST_HEADER_1~q ),
	.datab(\read_data_length[0]~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\read_data_length[0]~2_combout ),
	.cout());
defparam \read_data_length[0]~2 .lut_mask = 16'hEEEE;
defparam \read_data_length[0]~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \write_data_length[0]~0 (
	.dataa(\write_state.ST_HEADER_2~q ),
	.datab(\Add1~0_combout ),
	.datac(\header_in_bit_counter[2]~q ),
	.datad(\header_in_bit_counter[3]~q ),
	.cin(gnd),
	.combout(\write_data_length[0]~0_combout ),
	.cout());
defparam \write_data_length[0]~0 .lut_mask = 16'hEFFF;
defparam \write_data_length[0]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \write_state~17 (
	.dataa(\write_state~16_combout ),
	.datab(\read_data_length[0]~2_combout ),
	.datac(\write_data_length[0]~0_combout ),
	.datad(virtual_state_sdr),
	.cin(gnd),
	.combout(\write_state~17_combout ),
	.cout());
defparam \write_state~17 .lut_mask = 16'hFFBF;
defparam \write_state~17 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \write_state~20 (
	.dataa(\Equal6~2_combout ),
	.datab(\write_state~17_combout ),
	.datac(gnd),
	.datad(\write_state.ST_BYPASS~q ),
	.cin(gnd),
	.combout(\write_state~20_combout ),
	.cout());
defparam \write_state~20 .lut_mask = 16'h88BB;
defparam \write_state~20 .sum_lutc_input = "datac";

dffeas \write_state.ST_HEADER_1 (
	.clk(altera_internal_jtag),
	.d(\write_state~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_state~19_combout ),
	.q(\write_state.ST_HEADER_1~q ),
	.prn(vcc));
defparam \write_state.ST_HEADER_1 .is_wysiwyg = "true";
defparam \write_state.ST_HEADER_1 .power_up = "low";

fiftyfivenm_lcell_comb \read_data_length[0]~1 (
	.dataa(virtual_state_sdr),
	.datab(\Equal14~0_combout ),
	.datac(\write_state.ST_HEADER_1~q ),
	.datad(\read_data_length[0]~0_combout ),
	.cin(gnd),
	.combout(\read_data_length[0]~1_combout ),
	.cout());
defparam \read_data_length[0]~1 .lut_mask = 16'hFFFD;
defparam \read_data_length[0]~1 .sum_lutc_input = "datac";

dffeas \read_data_length[2] (
	.clk(altera_internal_jtag),
	.d(altera_internal_jtag1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\read_data_length[0]~1_combout ),
	.q(\read_data_length[2]~q ),
	.prn(vcc));
defparam \read_data_length[2] .is_wysiwyg = "true";
defparam \read_data_length[2] .power_up = "low";

fiftyfivenm_lcell_comb \header_in[14]~0 (
	.dataa(virtual_state_sdr),
	.datab(\Equal14~0_combout ),
	.datac(\write_state.ST_BYPASS~q ),
	.datad(\write_state.ST_WRITE_DATA~q ),
	.cin(gnd),
	.combout(\header_in[14]~0_combout ),
	.cout());
defparam \header_in[14]~0 .lut_mask = 16'hFDFF;
defparam \header_in[14]~0 .sum_lutc_input = "datac";

dffeas \header_in[15] (
	.clk(altera_internal_jtag),
	.d(altera_internal_jtag1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\header_in[14]~0_combout ),
	.q(\header_in[15]~q ),
	.prn(vcc));
defparam \header_in[15] .is_wysiwyg = "true";
defparam \header_in[15] .power_up = "low";

dffeas \header_in[14] (
	.clk(altera_internal_jtag),
	.d(\header_in[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\header_in[14]~0_combout ),
	.q(\header_in[14]~q ),
	.prn(vcc));
defparam \header_in[14] .is_wysiwyg = "true";
defparam \header_in[14] .power_up = "low";

dffeas \read_data_length[0] (
	.clk(altera_internal_jtag),
	.d(\header_in[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\read_data_length[0]~1_combout ),
	.q(\read_data_length[0]~q ),
	.prn(vcc));
defparam \read_data_length[0] .is_wysiwyg = "true";
defparam \read_data_length[0] .power_up = "low";

dffeas \read_data_length[1] (
	.clk(altera_internal_jtag),
	.d(\header_in[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\read_data_length[0]~1_combout ),
	.q(\read_data_length[1]~q ),
	.prn(vcc));
defparam \read_data_length[1] .is_wysiwyg = "true";
defparam \read_data_length[1] .power_up = "low";

fiftyfivenm_lcell_comb \read_data_all_valid~1 (
	.dataa(\read_data_length[2]~q ),
	.datab(\read_data_length[0]~q ),
	.datac(\read_data_length[1]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\read_data_all_valid~1_combout ),
	.cout());
defparam \read_data_all_valid~1 .lut_mask = 16'hFEFE;
defparam \read_data_all_valid~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \decode_header_1~2 (
	.dataa(virtual_state_cdr),
	.datab(\decode_header_1~q ),
	.datac(\write_state.ST_HEADER_1~q ),
	.datad(\header_in_bit_counter~2_combout ),
	.cin(gnd),
	.combout(\decode_header_1~2_combout ),
	.cout());
defparam \decode_header_1~2 .lut_mask = 16'hFEFF;
defparam \decode_header_1~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \decode_header_1~3 (
	.dataa(\write_state.ST_HEADER_1~q ),
	.datab(\read_data_length[0]~0_combout ),
	.datac(\decode_header_1~2_combout ),
	.datad(virtual_state_sdr),
	.cin(gnd),
	.combout(\decode_header_1~3_combout ),
	.cout());
defparam \decode_header_1~3 .lut_mask = 16'hFEFF;
defparam \decode_header_1~3 .sum_lutc_input = "datac";

dffeas decode_header_1(
	.clk(altera_internal_jtag),
	.d(\decode_header_1~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal14~0_combout ),
	.q(\decode_header_1~q ),
	.prn(vcc));
defparam decode_header_1.is_wysiwyg = "true";
defparam decode_header_1.power_up = "low";

fiftyfivenm_lcell_comb \read_data_all_valid~2 (
	.dataa(\decode_header_1~q ),
	.datab(\write_state.ST_HEADER_2~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\read_data_all_valid~2_combout ),
	.cout());
defparam \read_data_all_valid~2 .lut_mask = 16'hEEEE;
defparam \read_data_all_valid~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \read_data_all_valid~3 (
	.dataa(\read_data_all_valid~0_combout ),
	.datab(virtual_state_sdr),
	.datac(\read_data_all_valid~1_combout ),
	.datad(\read_data_all_valid~2_combout ),
	.cin(gnd),
	.combout(\read_data_all_valid~3_combout ),
	.cout());
defparam \read_data_all_valid~3 .lut_mask = 16'hFFFB;
defparam \read_data_all_valid~3 .sum_lutc_input = "datac";

dffeas read_data_all_valid(
	.clk(altera_internal_jtag),
	.d(\read_data_all_valid~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal14~0_combout ),
	.q(\read_data_all_valid~q ),
	.prn(vcc));
defparam read_data_all_valid.is_wysiwyg = "true";
defparam read_data_all_valid.power_up = "low";

fiftyfivenm_lcell_comb \Add8~0 (
	.dataa(\padded_bit_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add8~0_combout ),
	.cout(\Add8~1 ));
defparam \Add8~0 .lut_mask = 16'h55AA;
defparam \Add8~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \header_out_bit_counter~0 (
	.dataa(\header_out_bit_counter[0]~q ),
	.datab(\read_state.ST_HEADER~q ),
	.datac(gnd),
	.datad(virtual_state_sdr),
	.cin(gnd),
	.combout(\header_out_bit_counter~0_combout ),
	.cout());
defparam \header_out_bit_counter~0 .lut_mask = 16'h77FF;
defparam \header_out_bit_counter~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \header_out_bit_counter[0]~1 (
	.dataa(\Equal14~0_combout ),
	.datab(virtual_state_sdr),
	.datac(\read_state.ST_HEADER~q ),
	.datad(virtual_state_cdr),
	.cin(gnd),
	.combout(\header_out_bit_counter[0]~1_combout ),
	.cout());
defparam \header_out_bit_counter[0]~1 .lut_mask = 16'hBFFF;
defparam \header_out_bit_counter[0]~1 .sum_lutc_input = "datac";

dffeas \header_out_bit_counter[0] (
	.clk(altera_internal_jtag),
	.d(\header_out_bit_counter~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\header_out_bit_counter[0]~1_combout ),
	.q(\header_out_bit_counter[0]~q ),
	.prn(vcc));
defparam \header_out_bit_counter[0] .is_wysiwyg = "true";
defparam \header_out_bit_counter[0] .power_up = "low";

fiftyfivenm_lcell_comb \header_out_bit_counter~4 (
	.dataa(virtual_state_sdr),
	.datab(\header_out_bit_counter[0]~q ),
	.datac(\header_out_bit_counter[1]~q ),
	.datad(\read_state.ST_HEADER~q ),
	.cin(gnd),
	.combout(\header_out_bit_counter~4_combout ),
	.cout());
defparam \header_out_bit_counter~4 .lut_mask = 16'h7DFF;
defparam \header_out_bit_counter~4 .sum_lutc_input = "datac";

dffeas \header_out_bit_counter[1] (
	.clk(altera_internal_jtag),
	.d(\header_out_bit_counter~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\header_out_bit_counter[0]~1_combout ),
	.q(\header_out_bit_counter[1]~q ),
	.prn(vcc));
defparam \header_out_bit_counter[1] .is_wysiwyg = "true";
defparam \header_out_bit_counter[1] .power_up = "low";

fiftyfivenm_lcell_comb \Add6~0 (
	.dataa(gnd),
	.datab(\header_out_bit_counter[0]~q ),
	.datac(\header_out_bit_counter[1]~q ),
	.datad(\header_out_bit_counter[2]~q ),
	.cin(gnd),
	.combout(\Add6~0_combout ),
	.cout());
defparam \Add6~0 .lut_mask = 16'hC33C;
defparam \Add6~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \header_out_bit_counter~2 (
	.dataa(virtual_state_sdr),
	.datab(gnd),
	.datac(\read_state.ST_HEADER~q ),
	.datad(\Add6~0_combout ),
	.cin(gnd),
	.combout(\header_out_bit_counter~2_combout ),
	.cout());
defparam \header_out_bit_counter~2 .lut_mask = 16'h5FFF;
defparam \header_out_bit_counter~2 .sum_lutc_input = "datac";

dffeas \header_out_bit_counter[2] (
	.clk(altera_internal_jtag),
	.d(\header_out_bit_counter~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\header_out_bit_counter[0]~1_combout ),
	.q(\header_out_bit_counter[2]~q ),
	.prn(vcc));
defparam \header_out_bit_counter[2] .is_wysiwyg = "true";
defparam \header_out_bit_counter[2] .power_up = "low";

fiftyfivenm_lcell_comb \Add6~1 (
	.dataa(\header_out_bit_counter[2]~q ),
	.datab(\header_out_bit_counter[0]~q ),
	.datac(\header_out_bit_counter[1]~q ),
	.datad(\header_out_bit_counter[3]~q ),
	.cin(gnd),
	.combout(\Add6~1_combout ),
	.cout());
defparam \Add6~1 .lut_mask = 16'h6996;
defparam \Add6~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \header_out_bit_counter~3 (
	.dataa(virtual_state_sdr),
	.datab(gnd),
	.datac(\read_state.ST_HEADER~q ),
	.datad(\Add6~1_combout ),
	.cin(gnd),
	.combout(\header_out_bit_counter~3_combout ),
	.cout());
defparam \header_out_bit_counter~3 .lut_mask = 16'h5FFF;
defparam \header_out_bit_counter~3 .sum_lutc_input = "datac";

dffeas \header_out_bit_counter[3] (
	.clk(altera_internal_jtag),
	.d(\header_out_bit_counter~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\header_out_bit_counter[0]~1_combout ),
	.q(\header_out_bit_counter[3]~q ),
	.prn(vcc));
defparam \header_out_bit_counter[3] .is_wysiwyg = "true";
defparam \header_out_bit_counter[3] .power_up = "low";

fiftyfivenm_lcell_comb \Equal16~0 (
	.dataa(\header_out_bit_counter[0]~q ),
	.datab(\header_out_bit_counter[2]~q ),
	.datac(\header_out_bit_counter[3]~q ),
	.datad(\header_out_bit_counter[1]~q ),
	.cin(gnd),
	.combout(\Equal16~0_combout ),
	.cout());
defparam \Equal16~0 .lut_mask = 16'hBFFF;
defparam \Equal16~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \read_state~11 (
	.dataa(\Equal16~0_combout ),
	.datab(virtual_state_cdr),
	.datac(virtual_state_sdr),
	.datad(\read_state.ST_HEADER~q ),
	.cin(gnd),
	.combout(\read_state~11_combout ),
	.cout());
defparam \read_state~11 .lut_mask = 16'hF7FF;
defparam \read_state~11 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \read_state~12 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(state_3),
	.datac(\read_state.ST_HEADER~q ),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\read_state~12_combout ),
	.cout());
defparam \read_state~12 .lut_mask = 16'hFEFF;
defparam \read_state~12 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dr_data_out[2]~18 (
	.dataa(\Equal16~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\read_state.ST_HEADER~q ),
	.cin(gnd),
	.combout(\dr_data_out[2]~18_combout ),
	.cout());
defparam \dr_data_out[2]~18 .lut_mask = 16'hAAFF;
defparam \dr_data_out[2]~18 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \read_state~14 (
	.dataa(virtual_state_sdr),
	.datab(\Equal17~0_combout ),
	.datac(\dr_data_out[2]~18_combout ),
	.datad(\read_state.ST_PADDED~q ),
	.cin(gnd),
	.combout(\read_state~14_combout ),
	.cout());
defparam \read_state~14 .lut_mask = 16'hFDFF;
defparam \read_state~14 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \read_state~9 (
	.dataa(\Equal17~0_combout ),
	.datab(\read_state.ST_PADDED~q ),
	.datac(\dr_data_out[2]~18_combout ),
	.datad(virtual_state_sdr),
	.cin(gnd),
	.combout(\read_state~9_combout ),
	.cout());
defparam \read_state~9 .lut_mask = 16'hFFBF;
defparam \read_state~9 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \read_state~10 (
	.dataa(virtual_state_cdr),
	.datab(\read_state~9_combout ),
	.datac(gnd),
	.datad(\Equal14~0_combout ),
	.cin(gnd),
	.combout(\read_state~10_combout ),
	.cout());
defparam \read_state~10 .lut_mask = 16'hFF77;
defparam \read_state~10 .sum_lutc_input = "datac";

dffeas \read_state.ST_PADDED (
	.clk(altera_internal_jtag),
	.d(\read_state~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\read_state~10_combout ),
	.q(\read_state.ST_PADDED~q ),
	.prn(vcc));
defparam \read_state.ST_PADDED .is_wysiwyg = "true";
defparam \read_state.ST_PADDED .power_up = "low";

fiftyfivenm_lcell_comb \read_state~8 (
	.dataa(\Equal17~0_combout ),
	.datab(\read_state.ST_PADDED~q ),
	.datac(\dr_data_out[2]~18_combout ),
	.datad(virtual_state_sdr),
	.cin(gnd),
	.combout(\read_state~8_combout ),
	.cout());
defparam \read_state~8 .lut_mask = 16'hFDFF;
defparam \read_state~8 .sum_lutc_input = "datac";

dffeas \read_state.ST_READ_DATA (
	.clk(altera_internal_jtag),
	.d(\read_state~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\read_state~10_combout ),
	.q(\read_state.ST_READ_DATA~q ),
	.prn(vcc));
defparam \read_state.ST_READ_DATA .is_wysiwyg = "true";
defparam \read_state.ST_READ_DATA .power_up = "low";

fiftyfivenm_lcell_comb \read_state~13 (
	.dataa(\read_state~11_combout ),
	.datab(\read_state~12_combout ),
	.datac(\Equal17~0_combout ),
	.datad(\read_state.ST_READ_DATA~q ),
	.cin(gnd),
	.combout(\read_state~13_combout ),
	.cout());
defparam \read_state~13 .lut_mask = 16'h7FFF;
defparam \read_state~13 .sum_lutc_input = "datac";

dffeas \read_state.ST_HEADER (
	.clk(altera_internal_jtag),
	.d(\read_state~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal14~0_combout ),
	.q(\read_state.ST_HEADER~q ),
	.prn(vcc));
defparam \read_state.ST_HEADER .is_wysiwyg = "true";
defparam \read_state.ST_HEADER .power_up = "low";

fiftyfivenm_lcell_comb \padded_bit_counter[0]~0 (
	.dataa(virtual_state_sdr),
	.datab(\read_state.ST_HEADER~q ),
	.datac(\Equal17~0_combout ),
	.datad(\Equal16~0_combout ),
	.cin(gnd),
	.combout(\padded_bit_counter[0]~0_combout ),
	.cout());
defparam \padded_bit_counter[0]~0 .lut_mask = 16'hFFFD;
defparam \padded_bit_counter[0]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \padded_bit_counter~1 (
	.dataa(\Add8~0_combout ),
	.datab(\padded_bit_counter[0]~0_combout ),
	.datac(gnd),
	.datad(\read_state.ST_READ_DATA~q ),
	.cin(gnd),
	.combout(\padded_bit_counter~1_combout ),
	.cout());
defparam \padded_bit_counter~1 .lut_mask = 16'hEEFF;
defparam \padded_bit_counter~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \padded_bit_counter[0]~2 (
	.dataa(\Equal14~0_combout ),
	.datab(\padded_bit_counter[0]~0_combout ),
	.datac(\read_state.ST_READ_DATA~q ),
	.datad(virtual_state_cdr),
	.cin(gnd),
	.combout(\padded_bit_counter[0]~2_combout ),
	.cout());
defparam \padded_bit_counter[0]~2 .lut_mask = 16'hEFFF;
defparam \padded_bit_counter[0]~2 .sum_lutc_input = "datac";

dffeas \padded_bit_counter[0] (
	.clk(altera_internal_jtag),
	.d(\padded_bit_counter~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\padded_bit_counter[0]~2_combout ),
	.q(\padded_bit_counter[0]~q ),
	.prn(vcc));
defparam \padded_bit_counter[0] .is_wysiwyg = "true";
defparam \padded_bit_counter[0] .power_up = "low";

fiftyfivenm_lcell_comb \Add8~2 (
	.dataa(\padded_bit_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add8~1 ),
	.combout(\Add8~2_combout ),
	.cout(\Add8~3 ));
defparam \Add8~2 .lut_mask = 16'h5A5F;
defparam \Add8~2 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \padded_bit_counter~3 (
	.dataa(\padded_bit_counter[0]~0_combout ),
	.datab(\Add8~2_combout ),
	.datac(gnd),
	.datad(\read_state.ST_READ_DATA~q ),
	.cin(gnd),
	.combout(\padded_bit_counter~3_combout ),
	.cout());
defparam \padded_bit_counter~3 .lut_mask = 16'hEEFF;
defparam \padded_bit_counter~3 .sum_lutc_input = "datac";

dffeas \padded_bit_counter[1] (
	.clk(altera_internal_jtag),
	.d(\padded_bit_counter~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\padded_bit_counter[0]~2_combout ),
	.q(\padded_bit_counter[1]~q ),
	.prn(vcc));
defparam \padded_bit_counter[1] .is_wysiwyg = "true";
defparam \padded_bit_counter[1] .power_up = "low";

fiftyfivenm_lcell_comb \Add8~4 (
	.dataa(\padded_bit_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add8~3 ),
	.combout(\Add8~4_combout ),
	.cout(\Add8~5 ));
defparam \Add8~4 .lut_mask = 16'h5AAF;
defparam \Add8~4 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \padded_bit_counter~4 (
	.dataa(\padded_bit_counter[0]~0_combout ),
	.datab(\Add8~4_combout ),
	.datac(gnd),
	.datad(\read_state.ST_READ_DATA~q ),
	.cin(gnd),
	.combout(\padded_bit_counter~4_combout ),
	.cout());
defparam \padded_bit_counter~4 .lut_mask = 16'hEEFF;
defparam \padded_bit_counter~4 .sum_lutc_input = "datac";

dffeas \padded_bit_counter[2] (
	.clk(altera_internal_jtag),
	.d(\padded_bit_counter~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\padded_bit_counter[0]~2_combout ),
	.q(\padded_bit_counter[2]~q ),
	.prn(vcc));
defparam \padded_bit_counter[2] .is_wysiwyg = "true";
defparam \padded_bit_counter[2] .power_up = "low";

fiftyfivenm_lcell_comb \Add5~0 (
	.dataa(\offset[3]~q ),
	.datab(\Equal6~0_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add5~0_combout ),
	.cout(\Add5~1 ));
defparam \Add5~0 .lut_mask = 16'h66BB;
defparam \Add5~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add8~6 (
	.dataa(\padded_bit_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add8~5 ),
	.combout(\Add8~6_combout ),
	.cout(\Add8~7 ));
defparam \Add8~6 .lut_mask = 16'h5A5F;
defparam \Add8~6 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \padded_bit_counter~5 (
	.dataa(\Add5~0_combout ),
	.datab(\Add8~6_combout ),
	.datac(\padded_bit_counter[0]~0_combout ),
	.datad(\read_state.ST_READ_DATA~q ),
	.cin(gnd),
	.combout(\padded_bit_counter~5_combout ),
	.cout());
defparam \padded_bit_counter~5 .lut_mask = 16'hEFFE;
defparam \padded_bit_counter~5 .sum_lutc_input = "datac";

dffeas \padded_bit_counter[3] (
	.clk(altera_internal_jtag),
	.d(\padded_bit_counter~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\padded_bit_counter[0]~2_combout ),
	.q(\padded_bit_counter[3]~q ),
	.prn(vcc));
defparam \padded_bit_counter[3] .is_wysiwyg = "true";
defparam \padded_bit_counter[3] .power_up = "low";

fiftyfivenm_lcell_comb \Add5~2 (
	.dataa(\offset[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add5~1 ),
	.combout(\Add5~2_combout ),
	.cout(\Add5~3 ));
defparam \Add5~2 .lut_mask = 16'h5A5F;
defparam \Add5~2 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add8~8 (
	.dataa(\padded_bit_counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add8~7 ),
	.combout(\Add8~8_combout ),
	.cout(\Add8~9 ));
defparam \Add8~8 .lut_mask = 16'h5AAF;
defparam \Add8~8 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \padded_bit_counter~6 (
	.dataa(\Add5~2_combout ),
	.datab(\Add8~8_combout ),
	.datac(\padded_bit_counter[0]~0_combout ),
	.datad(\read_state.ST_READ_DATA~q ),
	.cin(gnd),
	.combout(\padded_bit_counter~6_combout ),
	.cout());
defparam \padded_bit_counter~6 .lut_mask = 16'hEFFE;
defparam \padded_bit_counter~6 .sum_lutc_input = "datac";

dffeas \padded_bit_counter[4] (
	.clk(altera_internal_jtag),
	.d(\padded_bit_counter~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\padded_bit_counter[0]~2_combout ),
	.q(\padded_bit_counter[4]~q ),
	.prn(vcc));
defparam \padded_bit_counter[4] .is_wysiwyg = "true";
defparam \padded_bit_counter[4] .power_up = "low";

fiftyfivenm_lcell_comb \idle_inserter_source_ready~0 (
	.dataa(\padded_bit_counter[1]~q ),
	.datab(\padded_bit_counter[2]~q ),
	.datac(\padded_bit_counter[3]~q ),
	.datad(\padded_bit_counter[4]~q ),
	.cin(gnd),
	.combout(\idle_inserter_source_ready~0_combout ),
	.cout());
defparam \idle_inserter_source_ready~0 .lut_mask = 16'h7FFF;
defparam \idle_inserter_source_ready~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add5~4 (
	.dataa(\offset[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add5~3 ),
	.combout(\Add5~4_combout ),
	.cout(\Add5~5 ));
defparam \Add5~4 .lut_mask = 16'h5AAF;
defparam \Add5~4 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add8~10 (
	.dataa(\padded_bit_counter[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add8~9 ),
	.combout(\Add8~10_combout ),
	.cout(\Add8~11 ));
defparam \Add8~10 .lut_mask = 16'h5A5F;
defparam \Add8~10 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \padded_bit_counter~7 (
	.dataa(\Add5~4_combout ),
	.datab(\Add8~10_combout ),
	.datac(\padded_bit_counter[0]~0_combout ),
	.datad(\read_state.ST_READ_DATA~q ),
	.cin(gnd),
	.combout(\padded_bit_counter~7_combout ),
	.cout());
defparam \padded_bit_counter~7 .lut_mask = 16'hEFFE;
defparam \padded_bit_counter~7 .sum_lutc_input = "datac";

dffeas \padded_bit_counter[5] (
	.clk(altera_internal_jtag),
	.d(\padded_bit_counter~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\padded_bit_counter[0]~2_combout ),
	.q(\padded_bit_counter[5]~q ),
	.prn(vcc));
defparam \padded_bit_counter[5] .is_wysiwyg = "true";
defparam \padded_bit_counter[5] .power_up = "low";

fiftyfivenm_lcell_comb \Add5~6 (
	.dataa(\offset[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add5~5 ),
	.combout(\Add5~6_combout ),
	.cout(\Add5~7 ));
defparam \Add5~6 .lut_mask = 16'h5A5F;
defparam \Add5~6 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add8~12 (
	.dataa(\padded_bit_counter[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add8~11 ),
	.combout(\Add8~12_combout ),
	.cout(\Add8~13 ));
defparam \Add8~12 .lut_mask = 16'h5AAF;
defparam \Add8~12 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \padded_bit_counter~8 (
	.dataa(\Add5~6_combout ),
	.datab(\Add8~12_combout ),
	.datac(\padded_bit_counter[0]~0_combout ),
	.datad(\read_state.ST_READ_DATA~q ),
	.cin(gnd),
	.combout(\padded_bit_counter~8_combout ),
	.cout());
defparam \padded_bit_counter~8 .lut_mask = 16'hEFFE;
defparam \padded_bit_counter~8 .sum_lutc_input = "datac";

dffeas \padded_bit_counter[6] (
	.clk(altera_internal_jtag),
	.d(\padded_bit_counter~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\padded_bit_counter[0]~2_combout ),
	.q(\padded_bit_counter[6]~q ),
	.prn(vcc));
defparam \padded_bit_counter[6] .is_wysiwyg = "true";
defparam \padded_bit_counter[6] .power_up = "low";

fiftyfivenm_lcell_comb \Add5~8 (
	.dataa(\offset[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add5~7 ),
	.combout(\Add5~8_combout ),
	.cout(\Add5~9 ));
defparam \Add5~8 .lut_mask = 16'h5AAF;
defparam \Add5~8 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add8~14 (
	.dataa(\padded_bit_counter[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add8~13 ),
	.combout(\Add8~14_combout ),
	.cout(\Add8~15 ));
defparam \Add8~14 .lut_mask = 16'h5A5F;
defparam \Add8~14 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \padded_bit_counter~9 (
	.dataa(\Add5~8_combout ),
	.datab(\Add8~14_combout ),
	.datac(\padded_bit_counter[0]~0_combout ),
	.datad(\read_state.ST_READ_DATA~q ),
	.cin(gnd),
	.combout(\padded_bit_counter~9_combout ),
	.cout());
defparam \padded_bit_counter~9 .lut_mask = 16'hEFFE;
defparam \padded_bit_counter~9 .sum_lutc_input = "datac";

dffeas \padded_bit_counter[7] (
	.clk(altera_internal_jtag),
	.d(\padded_bit_counter~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\padded_bit_counter[0]~2_combout ),
	.q(\padded_bit_counter[7]~q ),
	.prn(vcc));
defparam \padded_bit_counter[7] .is_wysiwyg = "true";
defparam \padded_bit_counter[7] .power_up = "low";

fiftyfivenm_lcell_comb \Add5~10 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add5~9 ),
	.combout(\Add5~10_combout ),
	.cout());
defparam \Add5~10 .lut_mask = 16'hF0F0;
defparam \Add5~10 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \padded_bit_counter~10 (
	.dataa(\padded_bit_counter[8]~q ),
	.datab(\Add5~10_combout ),
	.datac(gnd),
	.datad(virtual_state_cdr),
	.cin(gnd),
	.combout(\padded_bit_counter~10_combout ),
	.cout());
defparam \padded_bit_counter~10 .lut_mask = 16'hAACC;
defparam \padded_bit_counter~10 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add8~16 (
	.dataa(\padded_bit_counter[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add8~15 ),
	.combout(\Add8~16_combout ),
	.cout());
defparam \Add8~16 .lut_mask = 16'h5A5A;
defparam \Add8~16 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \dr_data_out[2]~11 (
	.dataa(\read_state.ST_READ_DATA~q ),
	.datab(\read_state.ST_HEADER~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\dr_data_out[2]~11_combout ),
	.cout());
defparam \dr_data_out[2]~11 .lut_mask = 16'hEEEE;
defparam \dr_data_out[2]~11 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \padded_bit_counter~11 (
	.dataa(\padded_bit_counter~10_combout ),
	.datab(\Add8~16_combout ),
	.datac(\padded_bit_counter[0]~0_combout ),
	.datad(\dr_data_out[2]~11_combout ),
	.cin(gnd),
	.combout(\padded_bit_counter~11_combout ),
	.cout());
defparam \padded_bit_counter~11 .lut_mask = 16'hEFFE;
defparam \padded_bit_counter~11 .sum_lutc_input = "datac";

dffeas \padded_bit_counter[8] (
	.clk(altera_internal_jtag),
	.d(\padded_bit_counter~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal14~0_combout ),
	.q(\padded_bit_counter[8]~q ),
	.prn(vcc));
defparam \padded_bit_counter[8] .is_wysiwyg = "true";
defparam \padded_bit_counter[8] .power_up = "low";

fiftyfivenm_lcell_comb \idle_inserter_source_ready~1 (
	.dataa(\padded_bit_counter[5]~q ),
	.datab(\padded_bit_counter[6]~q ),
	.datac(\padded_bit_counter[7]~q ),
	.datad(\padded_bit_counter[8]~q ),
	.cin(gnd),
	.combout(\idle_inserter_source_ready~1_combout ),
	.cout());
defparam \idle_inserter_source_ready~1 .lut_mask = 16'h7FFF;
defparam \idle_inserter_source_ready~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Equal17~0 (
	.dataa(\padded_bit_counter[0]~q ),
	.datab(gnd),
	.datac(\idle_inserter_source_ready~0_combout ),
	.datad(\idle_inserter_source_ready~1_combout ),
	.cin(gnd),
	.combout(\Equal17~0_combout ),
	.cout());
defparam \Equal17~0 .lut_mask = 16'hAFFF;
defparam \Equal17~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dr_data_out~7 (
	.dataa(\read_data_all_valid~q ),
	.datab(full1),
	.datac(gnd),
	.datad(\Equal17~0_combout ),
	.cin(gnd),
	.combout(\dr_data_out~7_combout ),
	.cout());
defparam \dr_data_out~7 .lut_mask = 16'hEEFF;
defparam \dr_data_out~7 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \read_data_bit_counter~0 (
	.dataa(\read_data_bit_counter[0]~q ),
	.datab(gnd),
	.datac(virtual_state_sdr),
	.datad(\read_state.ST_READ_DATA~q ),
	.cin(gnd),
	.combout(\read_data_bit_counter~0_combout ),
	.cout());
defparam \read_data_bit_counter~0 .lut_mask = 16'hFF5F;
defparam \read_data_bit_counter~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \read_data_bit_counter[0]~1 (
	.dataa(\Equal14~0_combout ),
	.datab(virtual_state_sdr),
	.datac(\read_state.ST_READ_DATA~q ),
	.datad(virtual_state_cdr),
	.cin(gnd),
	.combout(\read_data_bit_counter[0]~1_combout ),
	.cout());
defparam \read_data_bit_counter[0]~1 .lut_mask = 16'hFBFF;
defparam \read_data_bit_counter[0]~1 .sum_lutc_input = "datac";

dffeas \read_data_bit_counter[0] (
	.clk(altera_internal_jtag),
	.d(\read_data_bit_counter~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\read_data_bit_counter[0]~1_combout ),
	.q(\read_data_bit_counter[0]~q ),
	.prn(vcc));
defparam \read_data_bit_counter[0] .is_wysiwyg = "true";
defparam \read_data_bit_counter[0] .power_up = "low";

fiftyfivenm_lcell_comb \read_data_bit_counter~2 (
	.dataa(\read_data_bit_counter[0]~q ),
	.datab(\read_data_bit_counter[1]~q ),
	.datac(virtual_state_sdr),
	.datad(\read_state.ST_READ_DATA~q ),
	.cin(gnd),
	.combout(\read_data_bit_counter~2_combout ),
	.cout());
defparam \read_data_bit_counter~2 .lut_mask = 16'hFF6F;
defparam \read_data_bit_counter~2 .sum_lutc_input = "datac";

dffeas \read_data_bit_counter[1] (
	.clk(altera_internal_jtag),
	.d(\read_data_bit_counter~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\read_data_bit_counter[0]~1_combout ),
	.q(\read_data_bit_counter[1]~q ),
	.prn(vcc));
defparam \read_data_bit_counter[1] .is_wysiwyg = "true";
defparam \read_data_bit_counter[1] .power_up = "low";

fiftyfivenm_lcell_comb \Add9~0 (
	.dataa(gnd),
	.datab(\read_data_bit_counter[0]~q ),
	.datac(\read_data_bit_counter[1]~q ),
	.datad(\read_data_bit_counter[2]~q ),
	.cin(gnd),
	.combout(\Add9~0_combout ),
	.cout());
defparam \Add9~0 .lut_mask = 16'hC33C;
defparam \Add9~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \read_data_bit_counter~3 (
	.dataa(\Add9~0_combout ),
	.datab(gnd),
	.datac(virtual_state_sdr),
	.datad(\read_state.ST_READ_DATA~q ),
	.cin(gnd),
	.combout(\read_data_bit_counter~3_combout ),
	.cout());
defparam \read_data_bit_counter~3 .lut_mask = 16'hFF5F;
defparam \read_data_bit_counter~3 .sum_lutc_input = "datac";

dffeas \read_data_bit_counter[2] (
	.clk(altera_internal_jtag),
	.d(\read_data_bit_counter~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\read_data_bit_counter[0]~1_combout ),
	.q(\read_data_bit_counter[2]~q ),
	.prn(vcc));
defparam \read_data_bit_counter[2] .is_wysiwyg = "true";
defparam \read_data_bit_counter[2] .power_up = "low";

fiftyfivenm_lcell_comb \Equal1~0 (
	.dataa(\read_data_bit_counter[0]~q ),
	.datab(gnd),
	.datac(\read_data_bit_counter[1]~q ),
	.datad(\read_data_bit_counter[2]~q ),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
defparam \Equal1~0 .lut_mask = 16'hAFFF;
defparam \Equal1~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dr_data_out[2]~12 (
	.dataa(\Equal16~0_combout ),
	.datab(gnd),
	.datac(\read_state.ST_HEADER~q ),
	.datad(\read_state.ST_READ_DATA~q ),
	.cin(gnd),
	.combout(\dr_data_out[2]~12_combout ),
	.cout());
defparam \dr_data_out[2]~12 .lut_mask = 16'hA0AF;
defparam \dr_data_out[2]~12 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dr_data_out[2]~13 (
	.dataa(\Equal1~0_combout ),
	.datab(\dr_data_out[2]~11_combout ),
	.datac(\dr_data_out[2]~12_combout ),
	.datad(\Equal17~0_combout ),
	.cin(gnd),
	.combout(\dr_data_out[2]~13_combout ),
	.cout());
defparam \dr_data_out[2]~13 .lut_mask = 16'hFEFF;
defparam \dr_data_out[2]~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add10~0 (
	.dataa(\scan_length_byte_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add10~0_combout ),
	.cout(\Add10~1 ));
defparam \Add10~0 .lut_mask = 16'h55AA;
defparam \Add10~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \scan_length_byte_counter[0]~21 (
	.dataa(\scan_length_byte_counter[0]~q ),
	.datab(\scan_length_byte_counter[0]~12_combout ),
	.datac(\Add10~0_combout ),
	.datad(\scan_length_byte_counter[1]~11_combout ),
	.cin(gnd),
	.combout(\scan_length_byte_counter[0]~21_combout ),
	.cout());
defparam \scan_length_byte_counter[0]~21 .lut_mask = 16'hFFB8;
defparam \scan_length_byte_counter[0]~21 .sum_lutc_input = "datac";

dffeas \scan_length_byte_counter[0] (
	.clk(altera_internal_jtag),
	.d(\scan_length_byte_counter[0]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\scan_length_byte_counter[0]~q ),
	.prn(vcc));
defparam \scan_length_byte_counter[0] .is_wysiwyg = "true";
defparam \scan_length_byte_counter[0] .power_up = "low";

fiftyfivenm_lcell_comb \Add10~2 (
	.dataa(\scan_length_byte_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add10~1 ),
	.combout(\Add10~2_combout ),
	.cout(\Add10~3 ));
defparam \Add10~2 .lut_mask = 16'h5A5F;
defparam \Add10~2 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \scan_length_byte_counter[1]~13 (
	.dataa(\scan_length_byte_counter[1]~q ),
	.datab(\scan_length_byte_counter[0]~12_combout ),
	.datac(\Add10~2_combout ),
	.datad(\scan_length_byte_counter[1]~11_combout ),
	.cin(gnd),
	.combout(\scan_length_byte_counter[1]~13_combout ),
	.cout());
defparam \scan_length_byte_counter[1]~13 .lut_mask = 16'hFFB8;
defparam \scan_length_byte_counter[1]~13 .sum_lutc_input = "datac";

dffeas \scan_length_byte_counter[1] (
	.clk(altera_internal_jtag),
	.d(\scan_length_byte_counter[1]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\scan_length_byte_counter[1]~q ),
	.prn(vcc));
defparam \scan_length_byte_counter[1] .is_wysiwyg = "true";
defparam \scan_length_byte_counter[1] .power_up = "low";

fiftyfivenm_lcell_comb \Add10~4 (
	.dataa(\scan_length_byte_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add10~3 ),
	.combout(\Add10~4_combout ),
	.cout(\Add10~5 ));
defparam \Add10~4 .lut_mask = 16'h5AAF;
defparam \Add10~4 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \scan_length_byte_counter[2]~14 (
	.dataa(\scan_length_byte_counter[2]~q ),
	.datab(\scan_length_byte_counter[0]~12_combout ),
	.datac(\Add10~4_combout ),
	.datad(\scan_length_byte_counter[1]~11_combout ),
	.cin(gnd),
	.combout(\scan_length_byte_counter[2]~14_combout ),
	.cout());
defparam \scan_length_byte_counter[2]~14 .lut_mask = 16'hFFB8;
defparam \scan_length_byte_counter[2]~14 .sum_lutc_input = "datac";

dffeas \scan_length_byte_counter[2] (
	.clk(altera_internal_jtag),
	.d(\scan_length_byte_counter[2]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\scan_length_byte_counter[2]~q ),
	.prn(vcc));
defparam \scan_length_byte_counter[2] .is_wysiwyg = "true";
defparam \scan_length_byte_counter[2] .power_up = "low";

fiftyfivenm_lcell_comb \Add10~6 (
	.dataa(\scan_length_byte_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add10~5 ),
	.combout(\Add10~6_combout ),
	.cout(\Add10~7 ));
defparam \Add10~6 .lut_mask = 16'h5A5F;
defparam \Add10~6 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \scan_length_byte_counter[3]~15 (
	.dataa(\scan_length_byte_counter[3]~q ),
	.datab(\scan_length_byte_counter[0]~12_combout ),
	.datac(\Add10~6_combout ),
	.datad(\scan_length_byte_counter[1]~11_combout ),
	.cin(gnd),
	.combout(\scan_length_byte_counter[3]~15_combout ),
	.cout());
defparam \scan_length_byte_counter[3]~15 .lut_mask = 16'hFFB8;
defparam \scan_length_byte_counter[3]~15 .sum_lutc_input = "datac";

dffeas \scan_length_byte_counter[3] (
	.clk(altera_internal_jtag),
	.d(\scan_length_byte_counter[3]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\scan_length_byte_counter[3]~q ),
	.prn(vcc));
defparam \scan_length_byte_counter[3] .is_wysiwyg = "true";
defparam \scan_length_byte_counter[3] .power_up = "low";

fiftyfivenm_lcell_comb \Add10~8 (
	.dataa(\scan_length_byte_counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add10~7 ),
	.combout(\Add10~8_combout ),
	.cout(\Add10~9 ));
defparam \Add10~8 .lut_mask = 16'h5AAF;
defparam \Add10~8 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \scan_length_byte_counter[4]~16 (
	.dataa(\scan_length_byte_counter[4]~q ),
	.datab(\scan_length_byte_counter[0]~12_combout ),
	.datac(\Add10~8_combout ),
	.datad(\scan_length_byte_counter[1]~11_combout ),
	.cin(gnd),
	.combout(\scan_length_byte_counter[4]~16_combout ),
	.cout());
defparam \scan_length_byte_counter[4]~16 .lut_mask = 16'hFFB8;
defparam \scan_length_byte_counter[4]~16 .sum_lutc_input = "datac";

dffeas \scan_length_byte_counter[4] (
	.clk(altera_internal_jtag),
	.d(\scan_length_byte_counter[4]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\scan_length_byte_counter[4]~q ),
	.prn(vcc));
defparam \scan_length_byte_counter[4] .is_wysiwyg = "true";
defparam \scan_length_byte_counter[4] .power_up = "low";

fiftyfivenm_lcell_comb \Equal3~1 (
	.dataa(\scan_length_byte_counter[1]~q ),
	.datab(\scan_length_byte_counter[2]~q ),
	.datac(\scan_length_byte_counter[3]~q ),
	.datad(\scan_length_byte_counter[4]~q ),
	.cin(gnd),
	.combout(\Equal3~1_combout ),
	.cout());
defparam \Equal3~1 .lut_mask = 16'h7FFF;
defparam \Equal3~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add10~10 (
	.dataa(\scan_length_byte_counter[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add10~9 ),
	.combout(\Add10~10_combout ),
	.cout(\Add10~11 ));
defparam \Add10~10 .lut_mask = 16'h5A5F;
defparam \Add10~10 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \scan_length_byte_counter[5]~17 (
	.dataa(\scan_length_byte_counter[5]~q ),
	.datab(\scan_length_byte_counter[0]~12_combout ),
	.datac(\Add10~10_combout ),
	.datad(\scan_length_byte_counter[1]~11_combout ),
	.cin(gnd),
	.combout(\scan_length_byte_counter[5]~17_combout ),
	.cout());
defparam \scan_length_byte_counter[5]~17 .lut_mask = 16'hFFB8;
defparam \scan_length_byte_counter[5]~17 .sum_lutc_input = "datac";

dffeas \scan_length_byte_counter[5] (
	.clk(altera_internal_jtag),
	.d(\scan_length_byte_counter[5]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\scan_length_byte_counter[5]~q ),
	.prn(vcc));
defparam \scan_length_byte_counter[5] .is_wysiwyg = "true";
defparam \scan_length_byte_counter[5] .power_up = "low";

fiftyfivenm_lcell_comb \Add10~12 (
	.dataa(\scan_length_byte_counter[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add10~11 ),
	.combout(\Add10~12_combout ),
	.cout(\Add10~13 ));
defparam \Add10~12 .lut_mask = 16'h5AAF;
defparam \Add10~12 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \scan_length_byte_counter[6]~18 (
	.dataa(\scan_length_byte_counter[6]~q ),
	.datab(\scan_length_byte_counter[0]~12_combout ),
	.datac(\Add10~12_combout ),
	.datad(\scan_length_byte_counter[1]~11_combout ),
	.cin(gnd),
	.combout(\scan_length_byte_counter[6]~18_combout ),
	.cout());
defparam \scan_length_byte_counter[6]~18 .lut_mask = 16'hFFB8;
defparam \scan_length_byte_counter[6]~18 .sum_lutc_input = "datac";

dffeas \scan_length_byte_counter[6] (
	.clk(altera_internal_jtag),
	.d(\scan_length_byte_counter[6]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\scan_length_byte_counter[6]~q ),
	.prn(vcc));
defparam \scan_length_byte_counter[6] .is_wysiwyg = "true";
defparam \scan_length_byte_counter[6] .power_up = "low";

fiftyfivenm_lcell_comb \Equal3~2 (
	.dataa(\Equal3~1_combout ),
	.datab(\scan_length_byte_counter[5]~q ),
	.datac(\scan_length_byte_counter[6]~q ),
	.datad(\scan_length_byte_counter[7]~q ),
	.cin(gnd),
	.combout(\Equal3~2_combout ),
	.cout());
defparam \Equal3~2 .lut_mask = 16'hBFFF;
defparam \Equal3~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Equal3~0 (
	.dataa(\scan_length_byte_counter[11]~q ),
	.datab(\scan_length_byte_counter[12]~q ),
	.datac(\scan_length_byte_counter[13]~q ),
	.datad(\scan_length_byte_counter[14]~q ),
	.cin(gnd),
	.combout(\Equal3~0_combout ),
	.cout());
defparam \Equal3~0 .lut_mask = 16'h7FFF;
defparam \Equal3~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add10~28 (
	.dataa(\scan_length_byte_counter[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add10~27 ),
	.combout(\Add10~28_combout ),
	.cout(\Add10~29 ));
defparam \Add10~28 .lut_mask = 16'h5AAF;
defparam \Add10~28 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add10~30 (
	.dataa(\scan_length_byte_counter[15]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add10~29 ),
	.combout(\Add10~30_combout ),
	.cout(\Add10~31 ));
defparam \Add10~30 .lut_mask = 16'h5A5F;
defparam \Add10~30 .sum_lutc_input = "cin";

dffeas \header_in[13] (
	.clk(altera_internal_jtag),
	.d(\header_in[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\header_in[14]~0_combout ),
	.q(\header_in[13]~q ),
	.prn(vcc));
defparam \header_in[13] .is_wysiwyg = "true";
defparam \header_in[13] .power_up = "low";

dffeas \header_in[12] (
	.clk(altera_internal_jtag),
	.d(\header_in[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\header_in[14]~0_combout ),
	.q(\header_in[12]~q ),
	.prn(vcc));
defparam \header_in[12] .is_wysiwyg = "true";
defparam \header_in[12] .power_up = "low";

dffeas \header_in[11] (
	.clk(altera_internal_jtag),
	.d(\header_in[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\header_in[14]~0_combout ),
	.q(\header_in[11]~q ),
	.prn(vcc));
defparam \header_in[11] .is_wysiwyg = "true";
defparam \header_in[11] .power_up = "low";

dffeas \scan_length[7] (
	.clk(altera_internal_jtag),
	.d(\header_in[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\read_data_length[0]~1_combout ),
	.q(\scan_length[7]~q ),
	.prn(vcc));
defparam \scan_length[7] .is_wysiwyg = "true";
defparam \scan_length[7] .power_up = "low";

fiftyfivenm_lcell_comb \scan_length_byte_counter[15]~7 (
	.dataa(\Add10~30_combout ),
	.datab(\scan_length[7]~q ),
	.datac(gnd),
	.datad(\scan_length_byte_counter[1]~11_combout ),
	.cin(gnd),
	.combout(\scan_length_byte_counter[15]~7_combout ),
	.cout());
defparam \scan_length_byte_counter[15]~7 .lut_mask = 16'hAACC;
defparam \scan_length_byte_counter[15]~7 .sum_lutc_input = "datac";

dffeas \scan_length_byte_counter[15] (
	.clk(altera_internal_jtag),
	.d(\scan_length_byte_counter[15]~7_combout ),
	.asdata(\scan_length_byte_counter[15]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\scan_length_byte_counter[0]~12_combout ),
	.ena(vcc),
	.q(\scan_length_byte_counter[15]~q ),
	.prn(vcc));
defparam \scan_length_byte_counter[15] .is_wysiwyg = "true";
defparam \scan_length_byte_counter[15] .power_up = "low";

fiftyfivenm_lcell_comb \Add10~32 (
	.dataa(\scan_length_byte_counter[16]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add10~31 ),
	.combout(\Add10~32_combout ),
	.cout(\Add10~33 ));
defparam \Add10~32 .lut_mask = 16'h5AAF;
defparam \Add10~32 .sum_lutc_input = "cin";

dffeas \scan_length[8] (
	.clk(altera_internal_jtag),
	.d(\header_in[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\read_data_length[0]~1_combout ),
	.q(\scan_length[8]~q ),
	.prn(vcc));
defparam \scan_length[8] .is_wysiwyg = "true";
defparam \scan_length[8] .power_up = "low";

fiftyfivenm_lcell_comb \scan_length_byte_counter[16]~8 (
	.dataa(\Add10~32_combout ),
	.datab(\scan_length[8]~q ),
	.datac(gnd),
	.datad(\scan_length_byte_counter[1]~11_combout ),
	.cin(gnd),
	.combout(\scan_length_byte_counter[16]~8_combout ),
	.cout());
defparam \scan_length_byte_counter[16]~8 .lut_mask = 16'hAACC;
defparam \scan_length_byte_counter[16]~8 .sum_lutc_input = "datac";

dffeas \scan_length_byte_counter[16] (
	.clk(altera_internal_jtag),
	.d(\scan_length_byte_counter[16]~8_combout ),
	.asdata(\scan_length_byte_counter[16]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\scan_length_byte_counter[0]~12_combout ),
	.ena(vcc),
	.q(\scan_length_byte_counter[16]~q ),
	.prn(vcc));
defparam \scan_length_byte_counter[16] .is_wysiwyg = "true";
defparam \scan_length_byte_counter[16] .power_up = "low";

fiftyfivenm_lcell_comb \Add10~34 (
	.dataa(\scan_length_byte_counter[17]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add10~33 ),
	.combout(\Add10~34_combout ),
	.cout(\Add10~35 ));
defparam \Add10~34 .lut_mask = 16'h5A5F;
defparam \Add10~34 .sum_lutc_input = "cin";

dffeas \scan_length[9] (
	.clk(altera_internal_jtag),
	.d(\header_in[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\read_data_length[0]~1_combout ),
	.q(\scan_length[9]~q ),
	.prn(vcc));
defparam \scan_length[9] .is_wysiwyg = "true";
defparam \scan_length[9] .power_up = "low";

fiftyfivenm_lcell_comb \scan_length_byte_counter[17]~9 (
	.dataa(\Add10~34_combout ),
	.datab(\scan_length[9]~q ),
	.datac(gnd),
	.datad(\scan_length_byte_counter[1]~11_combout ),
	.cin(gnd),
	.combout(\scan_length_byte_counter[17]~9_combout ),
	.cout());
defparam \scan_length_byte_counter[17]~9 .lut_mask = 16'hAACC;
defparam \scan_length_byte_counter[17]~9 .sum_lutc_input = "datac";

dffeas \scan_length_byte_counter[17] (
	.clk(altera_internal_jtag),
	.d(\scan_length_byte_counter[17]~9_combout ),
	.asdata(\scan_length_byte_counter[17]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\scan_length_byte_counter[0]~12_combout ),
	.ena(vcc),
	.q(\scan_length_byte_counter[17]~q ),
	.prn(vcc));
defparam \scan_length_byte_counter[17] .is_wysiwyg = "true";
defparam \scan_length_byte_counter[17] .power_up = "low";

fiftyfivenm_lcell_comb \Add10~36 (
	.dataa(\scan_length_byte_counter[18]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add10~35 ),
	.combout(\Add10~36_combout ),
	.cout());
defparam \Add10~36 .lut_mask = 16'h5A5A;
defparam \Add10~36 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \scan_length_byte_counter[18]~20 (
	.dataa(\scan_length_byte_counter[18]~q ),
	.datab(\Add10~36_combout ),
	.datac(\scan_length_byte_counter[0]~12_combout ),
	.datad(\scan_length_byte_counter[1]~11_combout ),
	.cin(gnd),
	.combout(\scan_length_byte_counter[18]~20_combout ),
	.cout());
defparam \scan_length_byte_counter[18]~20 .lut_mask = 16'hACFF;
defparam \scan_length_byte_counter[18]~20 .sum_lutc_input = "datac";

dffeas \scan_length_byte_counter[18] (
	.clk(altera_internal_jtag),
	.d(\scan_length_byte_counter[18]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\scan_length_byte_counter[18]~q ),
	.prn(vcc));
defparam \scan_length_byte_counter[18] .is_wysiwyg = "true";
defparam \scan_length_byte_counter[18] .power_up = "low";

fiftyfivenm_lcell_comb \Equal3~3 (
	.dataa(\scan_length_byte_counter[18]~q ),
	.datab(\scan_length_byte_counter[15]~q ),
	.datac(\scan_length_byte_counter[16]~q ),
	.datad(\scan_length_byte_counter[17]~q ),
	.cin(gnd),
	.combout(\Equal3~3_combout ),
	.cout());
defparam \Equal3~3 .lut_mask = 16'h7FFF;
defparam \Equal3~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Equal3~4 (
	.dataa(\scan_length_byte_counter[0]~q ),
	.datab(\scan_length_byte_counter[8]~q ),
	.datac(\scan_length_byte_counter[9]~q ),
	.datad(\scan_length_byte_counter[10]~q ),
	.cin(gnd),
	.combout(\Equal3~4_combout ),
	.cout());
defparam \Equal3~4 .lut_mask = 16'h7FFF;
defparam \Equal3~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \scan_length_byte_counter[1]~10 (
	.dataa(\Equal3~0_combout ),
	.datab(\Equal3~3_combout ),
	.datac(\Equal3~4_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\scan_length_byte_counter[1]~10_combout ),
	.cout());
defparam \scan_length_byte_counter[1]~10 .lut_mask = 16'hFEFE;
defparam \scan_length_byte_counter[1]~10 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \scan_length_byte_counter[1]~11 (
	.dataa(\read_state.ST_READ_DATA~q ),
	.datab(\Equal1~0_combout ),
	.datac(\Equal3~2_combout ),
	.datad(\scan_length_byte_counter[1]~10_combout ),
	.cin(gnd),
	.combout(\scan_length_byte_counter[1]~11_combout ),
	.cout());
defparam \scan_length_byte_counter[1]~11 .lut_mask = 16'hFFF7;
defparam \scan_length_byte_counter[1]~11 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \scan_length_byte_counter[0]~12 (
	.dataa(virtual_state_sdr),
	.datab(\Equal14~0_combout ),
	.datac(\read_data_all_valid~2_combout ),
	.datad(\scan_length_byte_counter[1]~11_combout ),
	.cin(gnd),
	.combout(\scan_length_byte_counter[0]~12_combout ),
	.cout());
defparam \scan_length_byte_counter[0]~12 .lut_mask = 16'hFFBF;
defparam \scan_length_byte_counter[0]~12 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add10~14 (
	.dataa(\scan_length_byte_counter[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add10~13 ),
	.combout(\Add10~14_combout ),
	.cout(\Add10~15 ));
defparam \Add10~14 .lut_mask = 16'h5A5F;
defparam \Add10~14 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \scan_length_byte_counter[7]~19 (
	.dataa(\scan_length_byte_counter[7]~q ),
	.datab(\scan_length_byte_counter[0]~12_combout ),
	.datac(\Add10~14_combout ),
	.datad(\scan_length_byte_counter[1]~11_combout ),
	.cin(gnd),
	.combout(\scan_length_byte_counter[7]~19_combout ),
	.cout());
defparam \scan_length_byte_counter[7]~19 .lut_mask = 16'hFFB8;
defparam \scan_length_byte_counter[7]~19 .sum_lutc_input = "datac";

dffeas \scan_length_byte_counter[7] (
	.clk(altera_internal_jtag),
	.d(\scan_length_byte_counter[7]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\scan_length_byte_counter[7]~q ),
	.prn(vcc));
defparam \scan_length_byte_counter[7] .is_wysiwyg = "true";
defparam \scan_length_byte_counter[7] .power_up = "low";

fiftyfivenm_lcell_comb \Add10~16 (
	.dataa(\scan_length_byte_counter[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add10~15 ),
	.combout(\Add10~16_combout ),
	.cout(\Add10~17 ));
defparam \Add10~16 .lut_mask = 16'h5AAF;
defparam \Add10~16 .sum_lutc_input = "cin";

dffeas \header_in[10] (
	.clk(altera_internal_jtag),
	.d(\header_in[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\header_in[14]~0_combout ),
	.q(\header_in[10]~q ),
	.prn(vcc));
defparam \header_in[10] .is_wysiwyg = "true";
defparam \header_in[10] .power_up = "low";

dffeas \header_in[9] (
	.clk(altera_internal_jtag),
	.d(\header_in[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\header_in[14]~0_combout ),
	.q(\header_in[9]~q ),
	.prn(vcc));
defparam \header_in[9] .is_wysiwyg = "true";
defparam \header_in[9] .power_up = "low";

dffeas \header_in[8] (
	.clk(altera_internal_jtag),
	.d(\header_in[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\header_in[14]~0_combout ),
	.q(\header_in[8]~q ),
	.prn(vcc));
defparam \header_in[8] .is_wysiwyg = "true";
defparam \header_in[8] .power_up = "low";

dffeas \header_in[7] (
	.clk(altera_internal_jtag),
	.d(\header_in[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\header_in[14]~0_combout ),
	.q(\header_in[7]~q ),
	.prn(vcc));
defparam \header_in[7] .is_wysiwyg = "true";
defparam \header_in[7] .power_up = "low";

dffeas \header_in[6] (
	.clk(altera_internal_jtag),
	.d(\header_in[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\header_in[14]~0_combout ),
	.q(\header_in[6]~q ),
	.prn(vcc));
defparam \header_in[6] .is_wysiwyg = "true";
defparam \header_in[6] .power_up = "low";

dffeas \header_in[5] (
	.clk(altera_internal_jtag),
	.d(\header_in[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\header_in[14]~0_combout ),
	.q(\header_in[5]~q ),
	.prn(vcc));
defparam \header_in[5] .is_wysiwyg = "true";
defparam \header_in[5] .power_up = "low";

dffeas \header_in[4] (
	.clk(altera_internal_jtag),
	.d(\header_in[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\header_in[14]~0_combout ),
	.q(\header_in[4]~q ),
	.prn(vcc));
defparam \header_in[4] .is_wysiwyg = "true";
defparam \header_in[4] .power_up = "low";

dffeas \scan_length[0] (
	.clk(altera_internal_jtag),
	.d(\header_in[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\read_data_length[0]~1_combout ),
	.q(\scan_length[0]~q ),
	.prn(vcc));
defparam \scan_length[0] .is_wysiwyg = "true";
defparam \scan_length[0] .power_up = "low";

fiftyfivenm_lcell_comb \scan_length_byte_counter[8]~0 (
	.dataa(\Add10~16_combout ),
	.datab(\scan_length[0]~q ),
	.datac(gnd),
	.datad(\scan_length_byte_counter[1]~11_combout ),
	.cin(gnd),
	.combout(\scan_length_byte_counter[8]~0_combout ),
	.cout());
defparam \scan_length_byte_counter[8]~0 .lut_mask = 16'hAACC;
defparam \scan_length_byte_counter[8]~0 .sum_lutc_input = "datac";

dffeas \scan_length_byte_counter[8] (
	.clk(altera_internal_jtag),
	.d(\scan_length_byte_counter[8]~0_combout ),
	.asdata(\scan_length_byte_counter[8]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\scan_length_byte_counter[0]~12_combout ),
	.ena(vcc),
	.q(\scan_length_byte_counter[8]~q ),
	.prn(vcc));
defparam \scan_length_byte_counter[8] .is_wysiwyg = "true";
defparam \scan_length_byte_counter[8] .power_up = "low";

fiftyfivenm_lcell_comb \Add10~18 (
	.dataa(\scan_length_byte_counter[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add10~17 ),
	.combout(\Add10~18_combout ),
	.cout(\Add10~19 ));
defparam \Add10~18 .lut_mask = 16'h5A5F;
defparam \Add10~18 .sum_lutc_input = "cin";

dffeas \scan_length[1] (
	.clk(altera_internal_jtag),
	.d(\header_in[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\read_data_length[0]~1_combout ),
	.q(\scan_length[1]~q ),
	.prn(vcc));
defparam \scan_length[1] .is_wysiwyg = "true";
defparam \scan_length[1] .power_up = "low";

fiftyfivenm_lcell_comb \scan_length_byte_counter[9]~1 (
	.dataa(\Add10~18_combout ),
	.datab(\scan_length[1]~q ),
	.datac(gnd),
	.datad(\scan_length_byte_counter[1]~11_combout ),
	.cin(gnd),
	.combout(\scan_length_byte_counter[9]~1_combout ),
	.cout());
defparam \scan_length_byte_counter[9]~1 .lut_mask = 16'hAACC;
defparam \scan_length_byte_counter[9]~1 .sum_lutc_input = "datac";

dffeas \scan_length_byte_counter[9] (
	.clk(altera_internal_jtag),
	.d(\scan_length_byte_counter[9]~1_combout ),
	.asdata(\scan_length_byte_counter[9]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\scan_length_byte_counter[0]~12_combout ),
	.ena(vcc),
	.q(\scan_length_byte_counter[9]~q ),
	.prn(vcc));
defparam \scan_length_byte_counter[9] .is_wysiwyg = "true";
defparam \scan_length_byte_counter[9] .power_up = "low";

fiftyfivenm_lcell_comb \Add10~20 (
	.dataa(\scan_length_byte_counter[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add10~19 ),
	.combout(\Add10~20_combout ),
	.cout(\Add10~21 ));
defparam \Add10~20 .lut_mask = 16'h5AAF;
defparam \Add10~20 .sum_lutc_input = "cin";

dffeas \scan_length[2] (
	.clk(altera_internal_jtag),
	.d(\header_in[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\read_data_length[0]~1_combout ),
	.q(\scan_length[2]~q ),
	.prn(vcc));
defparam \scan_length[2] .is_wysiwyg = "true";
defparam \scan_length[2] .power_up = "low";

fiftyfivenm_lcell_comb \scan_length_byte_counter[10]~2 (
	.dataa(\Add10~20_combout ),
	.datab(\scan_length[2]~q ),
	.datac(gnd),
	.datad(\scan_length_byte_counter[1]~11_combout ),
	.cin(gnd),
	.combout(\scan_length_byte_counter[10]~2_combout ),
	.cout());
defparam \scan_length_byte_counter[10]~2 .lut_mask = 16'hAACC;
defparam \scan_length_byte_counter[10]~2 .sum_lutc_input = "datac";

dffeas \scan_length_byte_counter[10] (
	.clk(altera_internal_jtag),
	.d(\scan_length_byte_counter[10]~2_combout ),
	.asdata(\scan_length_byte_counter[10]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\scan_length_byte_counter[0]~12_combout ),
	.ena(vcc),
	.q(\scan_length_byte_counter[10]~q ),
	.prn(vcc));
defparam \scan_length_byte_counter[10] .is_wysiwyg = "true";
defparam \scan_length_byte_counter[10] .power_up = "low";

fiftyfivenm_lcell_comb \Add10~22 (
	.dataa(\scan_length_byte_counter[11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add10~21 ),
	.combout(\Add10~22_combout ),
	.cout(\Add10~23 ));
defparam \Add10~22 .lut_mask = 16'h5A5F;
defparam \Add10~22 .sum_lutc_input = "cin";

dffeas \scan_length[3] (
	.clk(altera_internal_jtag),
	.d(\header_in[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\read_data_length[0]~1_combout ),
	.q(\scan_length[3]~q ),
	.prn(vcc));
defparam \scan_length[3] .is_wysiwyg = "true";
defparam \scan_length[3] .power_up = "low";

fiftyfivenm_lcell_comb \scan_length_byte_counter[11]~3 (
	.dataa(\Add10~22_combout ),
	.datab(\scan_length[3]~q ),
	.datac(gnd),
	.datad(\scan_length_byte_counter[1]~11_combout ),
	.cin(gnd),
	.combout(\scan_length_byte_counter[11]~3_combout ),
	.cout());
defparam \scan_length_byte_counter[11]~3 .lut_mask = 16'hAACC;
defparam \scan_length_byte_counter[11]~3 .sum_lutc_input = "datac";

dffeas \scan_length_byte_counter[11] (
	.clk(altera_internal_jtag),
	.d(\scan_length_byte_counter[11]~3_combout ),
	.asdata(\scan_length_byte_counter[11]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\scan_length_byte_counter[0]~12_combout ),
	.ena(vcc),
	.q(\scan_length_byte_counter[11]~q ),
	.prn(vcc));
defparam \scan_length_byte_counter[11] .is_wysiwyg = "true";
defparam \scan_length_byte_counter[11] .power_up = "low";

fiftyfivenm_lcell_comb \Add10~24 (
	.dataa(\scan_length_byte_counter[12]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add10~23 ),
	.combout(\Add10~24_combout ),
	.cout(\Add10~25 ));
defparam \Add10~24 .lut_mask = 16'h5AAF;
defparam \Add10~24 .sum_lutc_input = "cin";

dffeas \scan_length[4] (
	.clk(altera_internal_jtag),
	.d(\header_in[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\read_data_length[0]~1_combout ),
	.q(\scan_length[4]~q ),
	.prn(vcc));
defparam \scan_length[4] .is_wysiwyg = "true";
defparam \scan_length[4] .power_up = "low";

fiftyfivenm_lcell_comb \scan_length_byte_counter[12]~4 (
	.dataa(\Add10~24_combout ),
	.datab(\scan_length[4]~q ),
	.datac(gnd),
	.datad(\scan_length_byte_counter[1]~11_combout ),
	.cin(gnd),
	.combout(\scan_length_byte_counter[12]~4_combout ),
	.cout());
defparam \scan_length_byte_counter[12]~4 .lut_mask = 16'hAACC;
defparam \scan_length_byte_counter[12]~4 .sum_lutc_input = "datac";

dffeas \scan_length_byte_counter[12] (
	.clk(altera_internal_jtag),
	.d(\scan_length_byte_counter[12]~4_combout ),
	.asdata(\scan_length_byte_counter[12]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\scan_length_byte_counter[0]~12_combout ),
	.ena(vcc),
	.q(\scan_length_byte_counter[12]~q ),
	.prn(vcc));
defparam \scan_length_byte_counter[12] .is_wysiwyg = "true";
defparam \scan_length_byte_counter[12] .power_up = "low";

fiftyfivenm_lcell_comb \Add10~26 (
	.dataa(\scan_length_byte_counter[13]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add10~25 ),
	.combout(\Add10~26_combout ),
	.cout(\Add10~27 ));
defparam \Add10~26 .lut_mask = 16'h5A5F;
defparam \Add10~26 .sum_lutc_input = "cin";

dffeas \scan_length[5] (
	.clk(altera_internal_jtag),
	.d(\header_in[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\read_data_length[0]~1_combout ),
	.q(\scan_length[5]~q ),
	.prn(vcc));
defparam \scan_length[5] .is_wysiwyg = "true";
defparam \scan_length[5] .power_up = "low";

fiftyfivenm_lcell_comb \scan_length_byte_counter[13]~5 (
	.dataa(\Add10~26_combout ),
	.datab(\scan_length[5]~q ),
	.datac(gnd),
	.datad(\scan_length_byte_counter[1]~11_combout ),
	.cin(gnd),
	.combout(\scan_length_byte_counter[13]~5_combout ),
	.cout());
defparam \scan_length_byte_counter[13]~5 .lut_mask = 16'hAACC;
defparam \scan_length_byte_counter[13]~5 .sum_lutc_input = "datac";

dffeas \scan_length_byte_counter[13] (
	.clk(altera_internal_jtag),
	.d(\scan_length_byte_counter[13]~5_combout ),
	.asdata(\scan_length_byte_counter[13]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\scan_length_byte_counter[0]~12_combout ),
	.ena(vcc),
	.q(\scan_length_byte_counter[13]~q ),
	.prn(vcc));
defparam \scan_length_byte_counter[13] .is_wysiwyg = "true";
defparam \scan_length_byte_counter[13] .power_up = "low";

dffeas \scan_length[6] (
	.clk(altera_internal_jtag),
	.d(\header_in[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\read_data_length[0]~1_combout ),
	.q(\scan_length[6]~q ),
	.prn(vcc));
defparam \scan_length[6] .is_wysiwyg = "true";
defparam \scan_length[6] .power_up = "low";

fiftyfivenm_lcell_comb \scan_length_byte_counter[14]~6 (
	.dataa(\Add10~28_combout ),
	.datab(\scan_length[6]~q ),
	.datac(gnd),
	.datad(\scan_length_byte_counter[1]~11_combout ),
	.cin(gnd),
	.combout(\scan_length_byte_counter[14]~6_combout ),
	.cout());
defparam \scan_length_byte_counter[14]~6 .lut_mask = 16'hAACC;
defparam \scan_length_byte_counter[14]~6 .sum_lutc_input = "datac";

dffeas \scan_length_byte_counter[14] (
	.clk(altera_internal_jtag),
	.d(\scan_length_byte_counter[14]~6_combout ),
	.asdata(\scan_length_byte_counter[14]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\scan_length_byte_counter[0]~12_combout ),
	.ena(vcc),
	.q(\scan_length_byte_counter[14]~q ),
	.prn(vcc));
defparam \scan_length_byte_counter[14] .is_wysiwyg = "true";
defparam \scan_length_byte_counter[14] .power_up = "low";

fiftyfivenm_lcell_comb \decoded_read_data_length[13]~0 (
	.dataa(\read_data_length[0]~q ),
	.datab(gnd),
	.datac(\read_data_length[2]~q ),
	.datad(\read_data_length[1]~q ),
	.cin(gnd),
	.combout(\decoded_read_data_length[13]~0_combout ),
	.cout());
defparam \decoded_read_data_length[13]~0 .lut_mask = 16'hAFFF;
defparam \decoded_read_data_length[13]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \decoded_read_data_length[12]~1 (
	.dataa(\read_data_length[2]~q ),
	.datab(\read_data_length[0]~q ),
	.datac(gnd),
	.datad(\read_data_length[1]~q ),
	.cin(gnd),
	.combout(\decoded_read_data_length[12]~1_combout ),
	.cout());
defparam \decoded_read_data_length[12]~1 .lut_mask = 16'hEEFF;
defparam \decoded_read_data_length[12]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \decoded_read_data_length[11]~2 (
	.dataa(\read_data_length[0]~q ),
	.datab(\read_data_length[1]~q ),
	.datac(gnd),
	.datad(\read_data_length[2]~q ),
	.cin(gnd),
	.combout(\decoded_read_data_length[11]~2_combout ),
	.cout());
defparam \decoded_read_data_length[11]~2 .lut_mask = 16'hEEFF;
defparam \decoded_read_data_length[11]~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \decoded_read_data_length[10]~3 (
	.dataa(\read_data_length[0]~q ),
	.datab(\read_data_length[1]~q ),
	.datac(gnd),
	.datad(\read_data_length[2]~q ),
	.cin(gnd),
	.combout(\decoded_read_data_length[10]~3_combout ),
	.cout());
defparam \decoded_read_data_length[10]~3 .lut_mask = 16'hEEFF;
defparam \decoded_read_data_length[10]~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \decoded_read_data_length[9]~4 (
	.dataa(\read_data_length[2]~q ),
	.datab(\read_data_length[0]~q ),
	.datac(gnd),
	.datad(\read_data_length[1]~q ),
	.cin(gnd),
	.combout(\decoded_read_data_length[9]~4_combout ),
	.cout());
defparam \decoded_read_data_length[9]~4 .lut_mask = 16'hEEFF;
defparam \decoded_read_data_length[9]~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \decoded_read_data_length[8]~5 (
	.dataa(\read_data_length[0]~q ),
	.datab(gnd),
	.datac(\read_data_length[2]~q ),
	.datad(\read_data_length[1]~q ),
	.cin(gnd),
	.combout(\decoded_read_data_length[8]~5_combout ),
	.cout());
defparam \decoded_read_data_length[8]~5 .lut_mask = 16'hAFFF;
defparam \decoded_read_data_length[8]~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \LessThan0~1 (
	.dataa(\Equal3~2_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\LessThan0~1_cout ));
defparam \LessThan0~1 .lut_mask = 16'h0055;
defparam \LessThan0~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \LessThan0~3 (
	.dataa(\decoded_read_data_length[8]~5_combout ),
	.datab(\scan_length_byte_counter[8]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~1_cout ),
	.combout(),
	.cout(\LessThan0~3_cout ));
defparam \LessThan0~3 .lut_mask = 16'h00BF;
defparam \LessThan0~3 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan0~5 (
	.dataa(\decoded_read_data_length[9]~4_combout ),
	.datab(\scan_length_byte_counter[9]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~3_cout ),
	.combout(),
	.cout(\LessThan0~5_cout ));
defparam \LessThan0~5 .lut_mask = 16'h00EF;
defparam \LessThan0~5 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan0~7 (
	.dataa(\decoded_read_data_length[10]~3_combout ),
	.datab(\scan_length_byte_counter[10]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~5_cout ),
	.combout(),
	.cout(\LessThan0~7_cout ));
defparam \LessThan0~7 .lut_mask = 16'h00BF;
defparam \LessThan0~7 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan0~9 (
	.dataa(\decoded_read_data_length[11]~2_combout ),
	.datab(\scan_length_byte_counter[11]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~7_cout ),
	.combout(),
	.cout(\LessThan0~9_cout ));
defparam \LessThan0~9 .lut_mask = 16'h00EF;
defparam \LessThan0~9 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan0~11 (
	.dataa(\decoded_read_data_length[12]~1_combout ),
	.datab(\scan_length_byte_counter[12]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~9_cout ),
	.combout(),
	.cout(\LessThan0~11_cout ));
defparam \LessThan0~11 .lut_mask = 16'h00BF;
defparam \LessThan0~11 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan0~13 (
	.dataa(\decoded_read_data_length[13]~0_combout ),
	.datab(\scan_length_byte_counter[13]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~11_cout ),
	.combout(),
	.cout(\LessThan0~13_cout ));
defparam \LessThan0~13 .lut_mask = 16'h00EF;
defparam \LessThan0~13 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \LessThan0~14 (
	.dataa(\read_data_all_valid~1_combout ),
	.datab(\scan_length_byte_counter[14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(\LessThan0~13_cout ),
	.combout(\LessThan0~14_combout ),
	.cout());
defparam \LessThan0~14 .lut_mask = 16'hFDFD;
defparam \LessThan0~14 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \read_data_valid~0 (
	.dataa(\read_data_bit_counter[1]~q ),
	.datab(\read_data_bit_counter[2]~q ),
	.datac(\read_data_bit_counter[0]~q ),
	.datad(\read_state.ST_HEADER~q ),
	.cin(gnd),
	.combout(\read_data_valid~0_combout ),
	.cout());
defparam \read_data_valid~0 .lut_mask = 16'hEFFF;
defparam \read_data_valid~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \read_data_valid~1 (
	.dataa(\Equal17~0_combout ),
	.datab(\dr_data_out[2]~12_combout ),
	.datac(virtual_state_sdr),
	.datad(\read_data_valid~0_combout ),
	.cin(gnd),
	.combout(\read_data_valid~1_combout ),
	.cout());
defparam \read_data_valid~1 .lut_mask = 16'h47FF;
defparam \read_data_valid~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \read_data_valid~2 (
	.dataa(\read_data_valid~q ),
	.datab(virtual_state_cdr),
	.datac(\Equal3~3_combout ),
	.datad(\read_data_valid~1_combout ),
	.cin(gnd),
	.combout(\read_data_valid~2_combout ),
	.cout());
defparam \read_data_valid~2 .lut_mask = 16'hFAFC;
defparam \read_data_valid~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \read_data_valid~3 (
	.dataa(\read_data_all_valid~q ),
	.datab(\LessThan0~14_combout ),
	.datac(\read_data_valid~1_combout ),
	.datad(\read_data_valid~2_combout ),
	.cin(gnd),
	.combout(\read_data_valid~3_combout ),
	.cout());
defparam \read_data_valid~3 .lut_mask = 16'hBFB3;
defparam \read_data_valid~3 .sum_lutc_input = "datac";

dffeas read_data_valid(
	.clk(altera_internal_jtag),
	.d(\read_data_valid~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal14~0_combout ),
	.q(\read_data_valid~q ),
	.prn(vcc));
defparam read_data_valid.is_wysiwyg = "true";
defparam read_data_valid.power_up = "low";

fiftyfivenm_lcell_comb \Equal3~5 (
	.dataa(\Equal3~0_combout ),
	.datab(\Equal3~2_combout ),
	.datac(\Equal3~3_combout ),
	.datad(\Equal3~4_combout ),
	.cin(gnd),
	.combout(\Equal3~5_combout ),
	.cout());
defparam \Equal3~5 .lut_mask = 16'hFFFE;
defparam \Equal3~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dr_data_out[2]~14 (
	.dataa(\read_state.ST_READ_DATA~q ),
	.datab(\read_data_valid~q ),
	.datac(gnd),
	.datad(\Equal3~5_combout ),
	.cin(gnd),
	.combout(\dr_data_out[2]~14_combout ),
	.cout());
defparam \dr_data_out[2]~14 .lut_mask = 16'hEEFF;
defparam \dr_data_out[2]~14 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dr_data_out[2]~15 (
	.dataa(full1),
	.datab(\dr_data_out[2]~14_combout ),
	.datac(\read_data_all_valid~q ),
	.datad(\read_state.ST_READ_DATA~q ),
	.cin(gnd),
	.combout(\dr_data_out[2]~15_combout ),
	.cout());
defparam \dr_data_out[2]~15 .lut_mask = 16'hFEFF;
defparam \dr_data_out[2]~15 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dr_data_out~16 (
	.dataa(\dr_data_out[2]~13_combout ),
	.datab(data1_1),
	.datac(out_data),
	.datad(\dr_data_out[2]~15_combout ),
	.cin(gnd),
	.combout(\dr_data_out~16_combout ),
	.cout());
defparam \dr_data_out~16 .lut_mask = 16'hEFFF;
defparam \dr_data_out~16 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dr_data_out[2]~9 (
	.dataa(gnd),
	.datab(\padded_bit_counter[0]~q ),
	.datac(\padded_bit_counter[1]~q ),
	.datad(\padded_bit_counter[2]~q ),
	.cin(gnd),
	.combout(\dr_data_out[2]~9_combout ),
	.cout());
defparam \dr_data_out[2]~9 .lut_mask = 16'h3FFF;
defparam \dr_data_out[2]~9 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dr_data_out[2]~19 (
	.dataa(\Equal17~0_combout ),
	.datab(\dr_data_out[2]~18_combout ),
	.datac(\dr_data_out[2]~9_combout ),
	.datad(\read_state.ST_PADDED~q ),
	.cin(gnd),
	.combout(\dr_data_out[2]~19_combout ),
	.cout());
defparam \dr_data_out[2]~19 .lut_mask = 16'hFFFE;
defparam \dr_data_out[2]~19 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dr_data_out~39 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(state_4),
	.datac(virtual_ir_scan_reg),
	.datad(\dr_data_out[2]~19_combout ),
	.cin(gnd),
	.combout(\dr_data_out~39_combout ),
	.cout());
defparam \dr_data_out~39 .lut_mask = 16'hEFFF;
defparam \dr_data_out~39 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dr_data_out[7]~10 (
	.dataa(full1),
	.datab(\Equal1~0_combout ),
	.datac(\read_data_valid~q ),
	.datad(\Equal3~5_combout ),
	.cin(gnd),
	.combout(\dr_data_out[7]~10_combout ),
	.cout());
defparam \dr_data_out[7]~10 .lut_mask = 16'hFEFF;
defparam \dr_data_out[7]~10 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dr_data_out[7]~36 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(state_4),
	.datac(data1_7),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\dr_data_out[7]~36_combout ),
	.cout());
defparam \dr_data_out[7]~36 .lut_mask = 16'hFEFF;
defparam \dr_data_out[7]~36 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dr_data_out[7]~40 (
	.dataa(\Equal16~0_combout ),
	.datab(\read_state.ST_HEADER~q ),
	.datac(\dr_data_out~7_combout ),
	.datad(\read_state.ST_READ_DATA~q ),
	.cin(gnd),
	.combout(\dr_data_out[7]~40_combout ),
	.cout());
defparam \dr_data_out[7]~40 .lut_mask = 16'hB8FF;
defparam \dr_data_out[7]~40 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dr_data_out[7]~37 (
	.dataa(\dr_data_out[7]~36_combout ),
	.datab(\dr_data_out[7]~40_combout ),
	.datac(\dr_data_out[7]~10_combout ),
	.datad(\dr_data_out[2]~11_combout ),
	.cin(gnd),
	.combout(\dr_data_out[7]~37_combout ),
	.cout());
defparam \dr_data_out[7]~37 .lut_mask = 16'hFFFE;
defparam \dr_data_out[7]~37 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dr_data_out[0]~38 (
	.dataa(irf_reg_2_1),
	.datab(irf_reg_0_1),
	.datac(irf_reg_1_1),
	.datad(\dr_info[4]~2_combout ),
	.cin(gnd),
	.combout(\dr_data_out[0]~38_combout ),
	.cout());
defparam \dr_data_out[0]~38 .lut_mask = 16'hFF7F;
defparam \dr_data_out[0]~38 .sum_lutc_input = "datac";

dffeas \dr_data_out[7] (
	.clk(altera_internal_jtag),
	.d(\dr_data_out[7]~37_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dr_data_out[0]~38_combout ),
	.q(\dr_data_out[7]~q ),
	.prn(vcc));
defparam \dr_data_out[7] .is_wysiwyg = "true";
defparam \dr_data_out[7] .power_up = "low";

fiftyfivenm_lcell_comb \dr_data_out~34 (
	.dataa(data1_6),
	.datab(\dr_data_out[7]~q ),
	.datac(gnd),
	.datad(\dr_data_out[2]~13_combout ),
	.cin(gnd),
	.combout(\dr_data_out~34_combout ),
	.cout());
defparam \dr_data_out~34 .lut_mask = 16'hAACC;
defparam \dr_data_out~34 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dr_data_out~24 (
	.dataa(\dr_data_out[2]~15_combout ),
	.datab(out_data),
	.datac(\dr_data_out[2]~13_combout ),
	.datad(\dr_data_out[2]~19_combout ),
	.cin(gnd),
	.combout(\dr_data_out~24_combout ),
	.cout());
defparam \dr_data_out~24 .lut_mask = 16'hBFFF;
defparam \dr_data_out~24 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dr_data_out~35 (
	.dataa(virtual_state_sdr),
	.datab(\dr_data_out~34_combout ),
	.datac(gnd),
	.datad(\dr_data_out~24_combout ),
	.cin(gnd),
	.combout(\dr_data_out~35_combout ),
	.cout());
defparam \dr_data_out~35 .lut_mask = 16'hDDFF;
defparam \dr_data_out~35 .sum_lutc_input = "datac";

dffeas \dr_data_out[6] (
	.clk(altera_internal_jtag),
	.d(\dr_data_out~35_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dr_data_out[0]~38_combout ),
	.q(\dr_data_out[6]~q ),
	.prn(vcc));
defparam \dr_data_out[6] .is_wysiwyg = "true";
defparam \dr_data_out[6] .power_up = "low";

fiftyfivenm_lcell_comb \dr_data_out[5]~28 (
	.dataa(\dr_data_out[7]~10_combout ),
	.datab(\idle_inserter|out_data~4_combout ),
	.datac(\dr_data_out[6]~q ),
	.datad(\Equal1~0_combout ),
	.cin(gnd),
	.combout(\dr_data_out[5]~28_combout ),
	.cout());
defparam \dr_data_out[5]~28 .lut_mask = 16'hFEFF;
defparam \dr_data_out[5]~28 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dr_data_out[5]~29 (
	.dataa(\dr_data_out[6]~q ),
	.datab(\padded_bit_counter[0]~q ),
	.datac(\padded_bit_counter[1]~q ),
	.datad(\padded_bit_counter[2]~q ),
	.cin(gnd),
	.combout(\dr_data_out[5]~29_combout ),
	.cout());
defparam \dr_data_out[5]~29 .lut_mask = 16'hFFFE;
defparam \dr_data_out[5]~29 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dr_data_out[5]~30 (
	.dataa(\read_data_all_valid~q ),
	.datab(full1),
	.datac(\idle_inserter|out_data~4_combout ),
	.datad(\Equal17~0_combout ),
	.cin(gnd),
	.combout(\dr_data_out[5]~30_combout ),
	.cout());
defparam \dr_data_out[5]~30 .lut_mask = 16'hFEFF;
defparam \dr_data_out[5]~30 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dr_data_out[5]~31 (
	.dataa(\dr_data_out[5]~28_combout ),
	.datab(\dr_data_out[5]~29_combout ),
	.datac(\dr_data_out[5]~30_combout ),
	.datad(\read_state.ST_READ_DATA~q ),
	.cin(gnd),
	.combout(\dr_data_out[5]~31_combout ),
	.cout());
defparam \dr_data_out[5]~31 .lut_mask = 16'hFAFC;
defparam \dr_data_out[5]~31 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dr_data_out[5]~32 (
	.dataa(\dr_data_out~7_combout ),
	.datab(\idle_inserter|out_data~4_combout ),
	.datac(\dr_data_out[6]~q ),
	.datad(\Equal16~0_combout ),
	.cin(gnd),
	.combout(\dr_data_out[5]~32_combout ),
	.cout());
defparam \dr_data_out[5]~32 .lut_mask = 16'hFAFC;
defparam \dr_data_out[5]~32 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dr_data_out[5]~33 (
	.dataa(virtual_state_sdr),
	.datab(\dr_data_out[5]~31_combout ),
	.datac(\dr_data_out[5]~32_combout ),
	.datad(\read_state.ST_HEADER~q ),
	.cin(gnd),
	.combout(\dr_data_out[5]~33_combout ),
	.cout());
defparam \dr_data_out[5]~33 .lut_mask = 16'hDDF5;
defparam \dr_data_out[5]~33 .sum_lutc_input = "datac";

dffeas \dr_data_out[5] (
	.clk(altera_internal_jtag),
	.d(\dr_data_out[5]~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dr_data_out[0]~38_combout ),
	.q(\dr_data_out[5]~q ),
	.prn(vcc));
defparam \dr_data_out[5] .is_wysiwyg = "true";
defparam \dr_data_out[5] .power_up = "low";

fiftyfivenm_lcell_comb \dr_data_out~26 (
	.dataa(\dr_data_out[5]~q ),
	.datab(\dr_data_out[2]~13_combout ),
	.datac(data1_4),
	.datad(out_data),
	.cin(gnd),
	.combout(\dr_data_out~26_combout ),
	.cout());
defparam \dr_data_out~26 .lut_mask = 16'hB8FF;
defparam \dr_data_out~26 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dr_data_out~27 (
	.dataa(\dr_data_out~39_combout ),
	.datab(\dr_data_out[2]~13_combout ),
	.datac(\dr_data_out[2]~15_combout ),
	.datad(\dr_data_out~26_combout ),
	.cin(gnd),
	.combout(\dr_data_out~27_combout ),
	.cout());
defparam \dr_data_out~27 .lut_mask = 16'hFFFB;
defparam \dr_data_out~27 .sum_lutc_input = "datac";

dffeas \dr_data_out[4] (
	.clk(altera_internal_jtag),
	.d(\dr_data_out~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dr_data_out[0]~38_combout ),
	.q(\dr_data_out[4]~q ),
	.prn(vcc));
defparam \dr_data_out[4] .is_wysiwyg = "true";
defparam \dr_data_out[4] .power_up = "low";

fiftyfivenm_lcell_comb \dr_data_out~23 (
	.dataa(data1_3),
	.datab(\dr_data_out[4]~q ),
	.datac(gnd),
	.datad(\dr_data_out[2]~13_combout ),
	.cin(gnd),
	.combout(\dr_data_out~23_combout ),
	.cout());
defparam \dr_data_out~23 .lut_mask = 16'hAACC;
defparam \dr_data_out~23 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dr_data_out~25 (
	.dataa(virtual_state_sdr),
	.datab(\dr_data_out~23_combout ),
	.datac(gnd),
	.datad(\dr_data_out~24_combout ),
	.cin(gnd),
	.combout(\dr_data_out~25_combout ),
	.cout());
defparam \dr_data_out~25 .lut_mask = 16'hDDFF;
defparam \dr_data_out~25 .sum_lutc_input = "datac";

dffeas \dr_data_out[3] (
	.clk(altera_internal_jtag),
	.d(\dr_data_out~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dr_data_out[0]~38_combout ),
	.q(\dr_data_out[3]~q ),
	.prn(vcc));
defparam \dr_data_out[3] .is_wysiwyg = "true";
defparam \dr_data_out[3] .power_up = "low";

fiftyfivenm_lcell_comb \dr_data_out~21 (
	.dataa(\dr_data_out[3]~q ),
	.datab(\dr_data_out[2]~13_combout ),
	.datac(data1_2),
	.datad(out_data),
	.cin(gnd),
	.combout(\dr_data_out~21_combout ),
	.cout());
defparam \dr_data_out~21 .lut_mask = 16'hFFB8;
defparam \dr_data_out~21 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dr_data_out~22 (
	.dataa(\dr_data_out~39_combout ),
	.datab(\dr_data_out[2]~13_combout ),
	.datac(\dr_data_out[2]~15_combout ),
	.datad(\dr_data_out~21_combout ),
	.cin(gnd),
	.combout(\dr_data_out~22_combout ),
	.cout());
defparam \dr_data_out~22 .lut_mask = 16'hFFFB;
defparam \dr_data_out~22 .sum_lutc_input = "datac";

dffeas \dr_data_out[2] (
	.clk(altera_internal_jtag),
	.d(\dr_data_out~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dr_data_out[0]~38_combout ),
	.q(\dr_data_out[2]~q ),
	.prn(vcc));
defparam \dr_data_out[2] .is_wysiwyg = "true";
defparam \dr_data_out[2] .power_up = "low";

fiftyfivenm_lcell_comb \dr_data_out~17 (
	.dataa(\dr_data_out[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\dr_data_out[2]~13_combout ),
	.cin(gnd),
	.combout(\dr_data_out~17_combout ),
	.cout());
defparam \dr_data_out~17 .lut_mask = 16'hAAFF;
defparam \dr_data_out~17 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dr_data_out~20 (
	.dataa(virtual_state_sdr),
	.datab(\dr_data_out~16_combout ),
	.datac(\dr_data_out~17_combout ),
	.datad(\dr_data_out[2]~19_combout ),
	.cin(gnd),
	.combout(\dr_data_out~20_combout ),
	.cout());
defparam \dr_data_out~20 .lut_mask = 16'hFFFD;
defparam \dr_data_out~20 .sum_lutc_input = "datac";

dffeas \dr_data_out[1] (
	.clk(altera_internal_jtag),
	.d(\dr_data_out~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dr_data_out[0]~38_combout ),
	.q(\dr_data_out[1]~q ),
	.prn(vcc));
defparam \dr_data_out[1] .is_wysiwyg = "true";
defparam \dr_data_out[1] .power_up = "low";

fiftyfivenm_lcell_comb \dr_data_out~8 (
	.dataa(\idle_inserter|out_data~3_combout ),
	.datab(\dr_data_out~7_combout ),
	.datac(\dr_data_out[1]~q ),
	.datad(\Equal16~0_combout ),
	.cin(gnd),
	.combout(\dr_data_out~8_combout ),
	.cout());
defparam \dr_data_out~8 .lut_mask = 16'hFAFC;
defparam \dr_data_out~8 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector41~2 (
	.dataa(\dr_data_out[1]~q ),
	.datab(\read_state.ST_READ_DATA~q ),
	.datac(\dr_data_out[2]~9_combout ),
	.datad(\Equal1~0_combout ),
	.cin(gnd),
	.combout(\Selector41~2_combout ),
	.cout());
defparam \Selector41~2 .lut_mask = 16'h8BFF;
defparam \Selector41~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector41~3 (
	.dataa(\dr_data_out[7]~10_combout ),
	.datab(\read_state.ST_READ_DATA~q ),
	.datac(\dr_data_out~7_combout ),
	.datad(\Equal17~0_combout ),
	.cin(gnd),
	.combout(\Selector41~3_combout ),
	.cout());
defparam \Selector41~3 .lut_mask = 16'hB8FF;
defparam \Selector41~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Selector41~4 (
	.dataa(data1_0),
	.datab(out_data),
	.datac(\Selector41~2_combout ),
	.datad(\Selector41~3_combout ),
	.cin(gnd),
	.combout(\Selector41~4_combout ),
	.cout());
defparam \Selector41~4 .lut_mask = 16'hFFFE;
defparam \Selector41~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dr_data_out[0]~0 (
	.dataa(\dr_data_out~8_combout ),
	.datab(\Selector41~4_combout ),
	.datac(gnd),
	.datad(\read_state.ST_HEADER~q ),
	.cin(gnd),
	.combout(\dr_data_out[0]~0_combout ),
	.cout());
defparam \dr_data_out[0]~0 .lut_mask = 16'hAACC;
defparam \dr_data_out[0]~0 .sum_lutc_input = "datac";

dffeas \dr_data_out[0] (
	.clk(altera_internal_jtag),
	.d(\dr_data_out[0]~0_combout ),
	.asdata(full1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(virtual_state_sdr),
	.ena(\dr_data_out[0]~38_combout ),
	.q(\dr_data_out[0]~q ),
	.prn(vcc));
defparam \dr_data_out[0] .is_wysiwyg = "true";
defparam \dr_data_out[0] .power_up = "low";

fiftyfivenm_lcell_comb \Mux0~0 (
	.dataa(irf_reg_1_1),
	.datab(\dr_loopback~q ),
	.datac(irf_reg_0_1),
	.datad(\dr_data_out[0]~q ),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
defparam \Mux0~0 .lut_mask = 16'hFFDE;
defparam \Mux0~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Equal14~1 (
	.dataa(irf_reg_0_1),
	.datab(irf_reg_1_1),
	.datac(gnd),
	.datad(irf_reg_2_1),
	.cin(gnd),
	.combout(\Equal14~1_combout ),
	.cout());
defparam \Equal14~1 .lut_mask = 16'hEEFF;
defparam \Equal14~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dr_info[8]~11 (
	.dataa(\dr_info[8]~q ),
	.datab(virtual_state_cdr),
	.datac(\Equal14~1_combout ),
	.datad(virtual_state_sdr),
	.cin(gnd),
	.combout(\dr_info[8]~11_combout ),
	.cout());
defparam \dr_info[8]~11 .lut_mask = 16'hBFB3;
defparam \dr_info[8]~11 .sum_lutc_input = "datac";

dffeas \dr_info[8] (
	.clk(altera_internal_jtag),
	.d(\dr_info[8]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dr_info[8]~q ),
	.prn(vcc));
defparam \dr_info[8] .is_wysiwyg = "true";
defparam \dr_info[8] .power_up = "low";

fiftyfivenm_lcell_comb \dr_info~10 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(state_4),
	.datac(\dr_info[8]~q ),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\dr_info~10_combout ),
	.cout());
defparam \dr_info~10 .lut_mask = 16'hFEFF;
defparam \dr_info~10 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dr_info[0]~12 (
	.dataa(irf_reg_0_1),
	.datab(irf_reg_1_1),
	.datac(irf_reg_2_1),
	.datad(\dr_info[4]~2_combout ),
	.cin(gnd),
	.combout(\dr_info[0]~12_combout ),
	.cout());
defparam \dr_info[0]~12 .lut_mask = 16'hFFEF;
defparam \dr_info[0]~12 .sum_lutc_input = "datac";

dffeas \dr_info[7] (
	.clk(altera_internal_jtag),
	.d(\dr_info~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dr_info[0]~12_combout ),
	.q(\dr_info[7]~q ),
	.prn(vcc));
defparam \dr_info[7] .is_wysiwyg = "true";
defparam \dr_info[7] .power_up = "low";

fiftyfivenm_lcell_comb \dr_info~9 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(state_4),
	.datac(\dr_info[7]~q ),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\dr_info~9_combout ),
	.cout());
defparam \dr_info~9 .lut_mask = 16'hFEFF;
defparam \dr_info~9 .sum_lutc_input = "datac";

dffeas \dr_info[6] (
	.clk(altera_internal_jtag),
	.d(\dr_info~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dr_info[0]~12_combout ),
	.q(\dr_info[6]~q ),
	.prn(vcc));
defparam \dr_info[6] .is_wysiwyg = "true";
defparam \dr_info[6] .power_up = "low";

fiftyfivenm_lcell_comb \dr_info~8 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(state_4),
	.datac(\dr_info[6]~q ),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\dr_info~8_combout ),
	.cout());
defparam \dr_info~8 .lut_mask = 16'hFEFF;
defparam \dr_info~8 .sum_lutc_input = "datac";

dffeas \dr_info[5] (
	.clk(altera_internal_jtag),
	.d(\dr_info~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dr_info[0]~12_combout ),
	.q(\dr_info[5]~q ),
	.prn(vcc));
defparam \dr_info[5] .is_wysiwyg = "true";
defparam \dr_info[5] .power_up = "low";

fiftyfivenm_lcell_comb \dr_info~7 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(state_4),
	.datac(\dr_info[5]~q ),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\dr_info~7_combout ),
	.cout());
defparam \dr_info~7 .lut_mask = 16'hFEFF;
defparam \dr_info~7 .sum_lutc_input = "datac";

dffeas \dr_info[4] (
	.clk(altera_internal_jtag),
	.d(\dr_info~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dr_info[0]~12_combout ),
	.q(\dr_info[4]~q ),
	.prn(vcc));
defparam \dr_info[4] .is_wysiwyg = "true";
defparam \dr_info[4] .power_up = "low";

fiftyfivenm_lcell_comb \dr_info~6 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(state_4),
	.datac(\dr_info[4]~q ),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\dr_info~6_combout ),
	.cout());
defparam \dr_info~6 .lut_mask = 16'hFEFF;
defparam \dr_info~6 .sum_lutc_input = "datac";

dffeas \dr_info[3] (
	.clk(altera_internal_jtag),
	.d(\dr_info~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dr_info[0]~12_combout ),
	.q(\dr_info[3]~q ),
	.prn(vcc));
defparam \dr_info[3] .is_wysiwyg = "true";
defparam \dr_info[3] .power_up = "low";

fiftyfivenm_lcell_comb \dr_info~5 (
	.dataa(virtual_ir_scan_reg),
	.datab(\dr_info[3]~q ),
	.datac(splitter_nodes_receive_0_3),
	.datad(state_4),
	.cin(gnd),
	.combout(\dr_info~5_combout ),
	.cout());
defparam \dr_info~5 .lut_mask = 16'hEFFF;
defparam \dr_info~5 .sum_lutc_input = "datac";

dffeas \dr_info[2] (
	.clk(altera_internal_jtag),
	.d(\dr_info~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dr_info[0]~12_combout ),
	.q(\dr_info[2]~q ),
	.prn(vcc));
defparam \dr_info[2] .is_wysiwyg = "true";
defparam \dr_info[2] .power_up = "low";

fiftyfivenm_lcell_comb \dr_info~4 (
	.dataa(virtual_ir_scan_reg),
	.datab(\dr_info[2]~q ),
	.datac(splitter_nodes_receive_0_3),
	.datad(state_4),
	.cin(gnd),
	.combout(\dr_info~4_combout ),
	.cout());
defparam \dr_info~4 .lut_mask = 16'hEFFF;
defparam \dr_info~4 .sum_lutc_input = "datac";

dffeas \dr_info[1] (
	.clk(altera_internal_jtag),
	.d(\dr_info~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dr_info[0]~12_combout ),
	.q(\dr_info[1]~q ),
	.prn(vcc));
defparam \dr_info[1] .is_wysiwyg = "true";
defparam \dr_info[1] .power_up = "low";

fiftyfivenm_lcell_comb \dr_info~3 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(state_4),
	.datac(\dr_info[1]~q ),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\dr_info~3_combout ),
	.cout());
defparam \dr_info~3 .lut_mask = 16'hFEFF;
defparam \dr_info~3 .sum_lutc_input = "datac";

dffeas \dr_info[0] (
	.clk(altera_internal_jtag),
	.d(\dr_info~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dr_info[0]~12_combout ),
	.q(\dr_info[0]~q ),
	.prn(vcc));
defparam \dr_info[0] .is_wysiwyg = "true";
defparam \dr_info[0] .power_up = "low";

fiftyfivenm_lcell_comb \Mux0~1 (
	.dataa(\dr_debug[0]~q ),
	.datab(irf_reg_1_1),
	.datac(\Mux0~0_combout ),
	.datad(\dr_info[0]~q ),
	.cin(gnd),
	.combout(\Mux0~1_combout ),
	.cout());
defparam \Mux0~1 .lut_mask = 16'hFFBE;
defparam \Mux0~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \idle_inserter_source_ready~2 (
	.dataa(\read_data_bit_counter[1]~q ),
	.datab(\read_state.ST_HEADER~q ),
	.datac(\read_data_bit_counter[0]~q ),
	.datad(\read_data_bit_counter[2]~q ),
	.cin(gnd),
	.combout(\idle_inserter_source_ready~2_combout ),
	.cout());
defparam \idle_inserter_source_ready~2 .lut_mask = 16'hEFFF;
defparam \idle_inserter_source_ready~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \idle_inserter_source_ready~3 (
	.dataa(\header_out_bit_counter[1]~q ),
	.datab(\header_out_bit_counter[2]~q ),
	.datac(\header_out_bit_counter[3]~q ),
	.datad(\header_out_bit_counter[0]~q ),
	.cin(gnd),
	.combout(\idle_inserter_source_ready~3_combout ),
	.cout());
defparam \idle_inserter_source_ready~3 .lut_mask = 16'hBFFF;
defparam \idle_inserter_source_ready~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \idle_inserter_source_ready~4 (
	.dataa(\padded_bit_counter[0]~q ),
	.datab(\read_state.ST_READ_DATA~q ),
	.datac(\idle_inserter_source_ready~0_combout ),
	.datad(\idle_inserter_source_ready~1_combout ),
	.cin(gnd),
	.combout(\idle_inserter_source_ready~4_combout ),
	.cout());
defparam \idle_inserter_source_ready~4 .lut_mask = 16'hFFFB;
defparam \idle_inserter_source_ready~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \idle_inserter_source_ready~5 (
	.dataa(\read_state.ST_HEADER~q ),
	.datab(\idle_inserter_source_ready~3_combout ),
	.datac(\Equal17~0_combout ),
	.datad(\idle_inserter_source_ready~4_combout ),
	.cin(gnd),
	.combout(\idle_inserter_source_ready~5_combout ),
	.cout());
defparam \idle_inserter_source_ready~5 .lut_mask = 16'hDF8F;
defparam \idle_inserter_source_ready~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \idle_inserter_source_ready~6 (
	.dataa(\read_data_all_valid~q ),
	.datab(\dr_data_out[2]~14_combout ),
	.datac(\idle_inserter_source_ready~2_combout ),
	.datad(\idle_inserter_source_ready~5_combout ),
	.cin(gnd),
	.combout(\idle_inserter_source_ready~6_combout ),
	.cout());
defparam \idle_inserter_source_ready~6 .lut_mask = 16'hFFFE;
defparam \idle_inserter_source_ready~6 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \idle_inserter_source_ready~7 (
	.dataa(virtual_state_sdr),
	.datab(\Equal14~0_combout ),
	.datac(\idle_inserter_source_ready~6_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\idle_inserter_source_ready~7_combout ),
	.cout());
defparam \idle_inserter_source_ready~7 .lut_mask = 16'hFDFD;
defparam \idle_inserter_source_ready~7 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \dr_data_in[1]~0 (
	.dataa(virtual_state_sdr),
	.datab(\Equal14~0_combout ),
	.datac(\write_state.ST_WRITE_DATA~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\dr_data_in[1]~0_combout ),
	.cout());
defparam \dr_data_in[1]~0 .lut_mask = 16'hFDFD;
defparam \dr_data_in[1]~0 .sum_lutc_input = "datac";

dffeas \dr_data_in[7] (
	.clk(altera_internal_jtag),
	.d(altera_internal_jtag1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dr_data_in[1]~0_combout ),
	.q(\dr_data_in[7]~q ),
	.prn(vcc));
defparam \dr_data_in[7] .is_wysiwyg = "true";
defparam \dr_data_in[7] .power_up = "low";

dffeas \dr_data_in[6] (
	.clk(altera_internal_jtag),
	.d(\dr_data_in[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dr_data_in[1]~0_combout ),
	.q(\dr_data_in[6]~q ),
	.prn(vcc));
defparam \dr_data_in[6] .is_wysiwyg = "true";
defparam \dr_data_in[6] .power_up = "low";

dffeas \dr_data_in[5] (
	.clk(altera_internal_jtag),
	.d(\dr_data_in[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dr_data_in[1]~0_combout ),
	.q(\dr_data_in[5]~q ),
	.prn(vcc));
defparam \dr_data_in[5] .is_wysiwyg = "true";
defparam \dr_data_in[5] .power_up = "low";

dffeas \dr_data_in[4] (
	.clk(altera_internal_jtag),
	.d(\dr_data_in[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dr_data_in[1]~0_combout ),
	.q(\dr_data_in[4]~q ),
	.prn(vcc));
defparam \dr_data_in[4] .is_wysiwyg = "true";
defparam \dr_data_in[4] .power_up = "low";

fiftyfivenm_lcell_comb \Add4~0 (
	.dataa(\valid_write_data_length_byte_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add4~0_combout ),
	.cout(\Add4~1 ));
defparam \Add4~0 .lut_mask = 16'h55AA;
defparam \Add4~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \valid_write_data_length_byte_counter~0 (
	.dataa(virtual_state_sdr),
	.datab(\write_state.ST_WRITE_DATA~q ),
	.datac(\always2~0_combout ),
	.datad(\Add4~0_combout ),
	.cin(gnd),
	.combout(\valid_write_data_length_byte_counter~0_combout ),
	.cout());
defparam \valid_write_data_length_byte_counter~0 .lut_mask = 16'hFFFD;
defparam \valid_write_data_length_byte_counter~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \decode_header_2~0 (
	.dataa(\write_state.ST_HEADER_2~q ),
	.datab(\write_state.ST_HEADER_1~q ),
	.datac(virtual_state_sdr),
	.datad(\write_state.ST_BYPASS~q ),
	.cin(gnd),
	.combout(\decode_header_2~0_combout ),
	.cout());
defparam \decode_header_2~0 .lut_mask = 16'hFEFF;
defparam \decode_header_2~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \decode_header_2~1 (
	.dataa(\decode_header_2~q ),
	.datab(virtual_ir_scan_reg),
	.datac(splitter_nodes_receive_0_3),
	.datad(state_3),
	.cin(gnd),
	.combout(\decode_header_2~1_combout ),
	.cout());
defparam \decode_header_2~1 .lut_mask = 16'hEFFF;
defparam \decode_header_2~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \decode_header_2~2 (
	.dataa(virtual_state_sdr),
	.datab(\decode_header_2~0_combout ),
	.datac(\decode_header_2~1_combout ),
	.datad(\write_data_length[0]~0_combout ),
	.cin(gnd),
	.combout(\decode_header_2~2_combout ),
	.cout());
defparam \decode_header_2~2 .lut_mask = 16'hFFFD;
defparam \decode_header_2~2 .sum_lutc_input = "datac";

dffeas decode_header_2(
	.clk(altera_internal_jtag),
	.d(\decode_header_2~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Equal14~0_combout ),
	.q(\decode_header_2~q ),
	.prn(vcc));
defparam decode_header_2.is_wysiwyg = "true";
defparam decode_header_2.power_up = "low";

fiftyfivenm_lcell_comb \valid_write_data_length_byte_counter[5]~1 (
	.dataa(virtual_state_sdr),
	.datab(\write_state.ST_WRITE_DATA~q ),
	.datac(\always2~0_combout ),
	.datad(\decode_header_2~q ),
	.cin(gnd),
	.combout(\valid_write_data_length_byte_counter[5]~1_combout ),
	.cout());
defparam \valid_write_data_length_byte_counter[5]~1 .lut_mask = 16'hFFFD;
defparam \valid_write_data_length_byte_counter[5]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \valid_write_data_length_byte_counter[0]~2 (
	.dataa(\Equal14~0_combout ),
	.datab(\valid_write_data_length_byte_counter[5]~1_combout ),
	.datac(gnd),
	.datad(virtual_state_cdr),
	.cin(gnd),
	.combout(\valid_write_data_length_byte_counter[0]~2_combout ),
	.cout());
defparam \valid_write_data_length_byte_counter[0]~2 .lut_mask = 16'hEEFF;
defparam \valid_write_data_length_byte_counter[0]~2 .sum_lutc_input = "datac";

dffeas \valid_write_data_length_byte_counter[0] (
	.clk(altera_internal_jtag),
	.d(\valid_write_data_length_byte_counter~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\valid_write_data_length_byte_counter[0]~2_combout ),
	.q(\valid_write_data_length_byte_counter[0]~q ),
	.prn(vcc));
defparam \valid_write_data_length_byte_counter[0] .is_wysiwyg = "true";
defparam \valid_write_data_length_byte_counter[0] .power_up = "low";

fiftyfivenm_lcell_comb \Add4~2 (
	.dataa(\valid_write_data_length_byte_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add4~1 ),
	.combout(\Add4~2_combout ),
	.cout(\Add4~3 ));
defparam \Add4~2 .lut_mask = 16'h5A5F;
defparam \Add4~2 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \valid_write_data_length_byte_counter~3 (
	.dataa(virtual_state_sdr),
	.datab(\write_state.ST_WRITE_DATA~q ),
	.datac(\always2~0_combout ),
	.datad(\Add4~2_combout ),
	.cin(gnd),
	.combout(\valid_write_data_length_byte_counter~3_combout ),
	.cout());
defparam \valid_write_data_length_byte_counter~3 .lut_mask = 16'hFFFD;
defparam \valid_write_data_length_byte_counter~3 .sum_lutc_input = "datac";

dffeas \valid_write_data_length_byte_counter[1] (
	.clk(altera_internal_jtag),
	.d(\valid_write_data_length_byte_counter~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\valid_write_data_length_byte_counter[0]~2_combout ),
	.q(\valid_write_data_length_byte_counter[1]~q ),
	.prn(vcc));
defparam \valid_write_data_length_byte_counter[1] .is_wysiwyg = "true";
defparam \valid_write_data_length_byte_counter[1] .power_up = "low";

fiftyfivenm_lcell_comb \Add4~4 (
	.dataa(\valid_write_data_length_byte_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add4~3 ),
	.combout(\Add4~4_combout ),
	.cout(\Add4~5 ));
defparam \Add4~4 .lut_mask = 16'h5AAF;
defparam \Add4~4 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \valid_write_data_length_byte_counter~4 (
	.dataa(virtual_state_sdr),
	.datab(\write_state.ST_WRITE_DATA~q ),
	.datac(\always2~0_combout ),
	.datad(\Add4~4_combout ),
	.cin(gnd),
	.combout(\valid_write_data_length_byte_counter~4_combout ),
	.cout());
defparam \valid_write_data_length_byte_counter~4 .lut_mask = 16'hFFFD;
defparam \valid_write_data_length_byte_counter~4 .sum_lutc_input = "datac";

dffeas \valid_write_data_length_byte_counter[2] (
	.clk(altera_internal_jtag),
	.d(\valid_write_data_length_byte_counter~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\valid_write_data_length_byte_counter[0]~2_combout ),
	.q(\valid_write_data_length_byte_counter[2]~q ),
	.prn(vcc));
defparam \valid_write_data_length_byte_counter[2] .is_wysiwyg = "true";
defparam \valid_write_data_length_byte_counter[2] .power_up = "low";

fiftyfivenm_lcell_comb \Add4~6 (
	.dataa(\valid_write_data_length_byte_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add4~5 ),
	.combout(\Add4~6_combout ),
	.cout(\Add4~7 ));
defparam \Add4~6 .lut_mask = 16'h5A5F;
defparam \Add4~6 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \valid_write_data_length_byte_counter~5 (
	.dataa(virtual_state_sdr),
	.datab(\write_state.ST_WRITE_DATA~q ),
	.datac(\always2~0_combout ),
	.datad(\Add4~6_combout ),
	.cin(gnd),
	.combout(\valid_write_data_length_byte_counter~5_combout ),
	.cout());
defparam \valid_write_data_length_byte_counter~5 .lut_mask = 16'hFFFD;
defparam \valid_write_data_length_byte_counter~5 .sum_lutc_input = "datac";

dffeas \valid_write_data_length_byte_counter[3] (
	.clk(altera_internal_jtag),
	.d(\valid_write_data_length_byte_counter~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\valid_write_data_length_byte_counter[0]~2_combout ),
	.q(\valid_write_data_length_byte_counter[3]~q ),
	.prn(vcc));
defparam \valid_write_data_length_byte_counter[3] .is_wysiwyg = "true";
defparam \valid_write_data_length_byte_counter[3] .power_up = "low";

fiftyfivenm_lcell_comb \Equal13~0 (
	.dataa(\valid_write_data_length_byte_counter[0]~q ),
	.datab(\valid_write_data_length_byte_counter[1]~q ),
	.datac(\valid_write_data_length_byte_counter[2]~q ),
	.datad(\valid_write_data_length_byte_counter[3]~q ),
	.cin(gnd),
	.combout(\Equal13~0_combout ),
	.cout());
defparam \Equal13~0 .lut_mask = 16'h7FFF;
defparam \Equal13~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add4~8 (
	.dataa(\valid_write_data_length_byte_counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add4~7 ),
	.combout(\Add4~8_combout ),
	.cout(\Add4~9 ));
defparam \Add4~8 .lut_mask = 16'h5AAF;
defparam \Add4~8 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \valid_write_data_length_byte_counter~6 (
	.dataa(virtual_state_sdr),
	.datab(\write_state.ST_WRITE_DATA~q ),
	.datac(\always2~0_combout ),
	.datad(\Add4~8_combout ),
	.cin(gnd),
	.combout(\valid_write_data_length_byte_counter~6_combout ),
	.cout());
defparam \valid_write_data_length_byte_counter~6 .lut_mask = 16'hFFFD;
defparam \valid_write_data_length_byte_counter~6 .sum_lutc_input = "datac";

dffeas \valid_write_data_length_byte_counter[4] (
	.clk(altera_internal_jtag),
	.d(\valid_write_data_length_byte_counter~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\valid_write_data_length_byte_counter[0]~2_combout ),
	.q(\valid_write_data_length_byte_counter[4]~q ),
	.prn(vcc));
defparam \valid_write_data_length_byte_counter[4] .is_wysiwyg = "true";
defparam \valid_write_data_length_byte_counter[4] .power_up = "low";

fiftyfivenm_lcell_comb \Add4~10 (
	.dataa(\valid_write_data_length_byte_counter[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add4~9 ),
	.combout(\Add4~10_combout ),
	.cout(\Add4~11 ));
defparam \Add4~10 .lut_mask = 16'h5A5F;
defparam \Add4~10 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \valid_write_data_length_byte_counter~7 (
	.dataa(virtual_state_sdr),
	.datab(\write_state.ST_WRITE_DATA~q ),
	.datac(\always2~0_combout ),
	.datad(\Add4~10_combout ),
	.cin(gnd),
	.combout(\valid_write_data_length_byte_counter~7_combout ),
	.cout());
defparam \valid_write_data_length_byte_counter~7 .lut_mask = 16'hFFFD;
defparam \valid_write_data_length_byte_counter~7 .sum_lutc_input = "datac";

dffeas \valid_write_data_length_byte_counter[5] (
	.clk(altera_internal_jtag),
	.d(\valid_write_data_length_byte_counter~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\valid_write_data_length_byte_counter[0]~2_combout ),
	.q(\valid_write_data_length_byte_counter[5]~q ),
	.prn(vcc));
defparam \valid_write_data_length_byte_counter[5] .is_wysiwyg = "true";
defparam \valid_write_data_length_byte_counter[5] .power_up = "low";

fiftyfivenm_lcell_comb \Add4~12 (
	.dataa(\valid_write_data_length_byte_counter[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add4~11 ),
	.combout(\Add4~12_combout ),
	.cout(\Add4~13 ));
defparam \Add4~12 .lut_mask = 16'h5AAF;
defparam \Add4~12 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \valid_write_data_length_byte_counter~8 (
	.dataa(virtual_state_sdr),
	.datab(\write_state.ST_WRITE_DATA~q ),
	.datac(\always2~0_combout ),
	.datad(\Add4~12_combout ),
	.cin(gnd),
	.combout(\valid_write_data_length_byte_counter~8_combout ),
	.cout());
defparam \valid_write_data_length_byte_counter~8 .lut_mask = 16'hFFFD;
defparam \valid_write_data_length_byte_counter~8 .sum_lutc_input = "datac";

dffeas \valid_write_data_length_byte_counter[6] (
	.clk(altera_internal_jtag),
	.d(\valid_write_data_length_byte_counter~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\valid_write_data_length_byte_counter[0]~2_combout ),
	.q(\valid_write_data_length_byte_counter[6]~q ),
	.prn(vcc));
defparam \valid_write_data_length_byte_counter[6] .is_wysiwyg = "true";
defparam \valid_write_data_length_byte_counter[6] .power_up = "low";

fiftyfivenm_lcell_comb \Add4~14 (
	.dataa(\valid_write_data_length_byte_counter[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add4~13 ),
	.combout(\Add4~14_combout ),
	.cout(\Add4~15 ));
defparam \Add4~14 .lut_mask = 16'h5A5F;
defparam \Add4~14 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \valid_write_data_length_byte_counter~9 (
	.dataa(\always2~0_combout ),
	.datab(\valid_write_data_length_byte_counter[5]~1_combout ),
	.datac(\Add4~14_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\valid_write_data_length_byte_counter~9_combout ),
	.cout());
defparam \valid_write_data_length_byte_counter~9 .lut_mask = 16'hFEFE;
defparam \valid_write_data_length_byte_counter~9 .sum_lutc_input = "datac";

dffeas \valid_write_data_length_byte_counter[7] (
	.clk(altera_internal_jtag),
	.d(\valid_write_data_length_byte_counter~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\valid_write_data_length_byte_counter[0]~2_combout ),
	.q(\valid_write_data_length_byte_counter[7]~q ),
	.prn(vcc));
defparam \valid_write_data_length_byte_counter[7] .is_wysiwyg = "true";
defparam \valid_write_data_length_byte_counter[7] .power_up = "low";

fiftyfivenm_lcell_comb \Equal13~1 (
	.dataa(\valid_write_data_length_byte_counter[4]~q ),
	.datab(\valid_write_data_length_byte_counter[5]~q ),
	.datac(\valid_write_data_length_byte_counter[6]~q ),
	.datad(\valid_write_data_length_byte_counter[7]~q ),
	.cin(gnd),
	.combout(\Equal13~1_combout ),
	.cout());
defparam \Equal13~1 .lut_mask = 16'h7FFF;
defparam \Equal13~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \write_data_length[0]~1 (
	.dataa(virtual_state_sdr),
	.datab(\Equal14~0_combout ),
	.datac(\write_data_length[0]~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\write_data_length[0]~1_combout ),
	.cout());
defparam \write_data_length[0]~1 .lut_mask = 16'hFDFD;
defparam \write_data_length[0]~1 .sum_lutc_input = "datac";

dffeas \write_data_length[0] (
	.clk(altera_internal_jtag),
	.d(\header_in[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_data_length[0]~1_combout ),
	.q(\write_data_length[0]~q ),
	.prn(vcc));
defparam \write_data_length[0] .is_wysiwyg = "true";
defparam \write_data_length[0] .power_up = "low";

fiftyfivenm_lcell_comb \valid_write_data_length_byte_counter~10 (
	.dataa(\write_data_length[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\always2~0_combout ),
	.cin(gnd),
	.combout(\valid_write_data_length_byte_counter~10_combout ),
	.cout());
defparam \valid_write_data_length_byte_counter~10 .lut_mask = 16'hAAFF;
defparam \valid_write_data_length_byte_counter~10 .sum_lutc_input = "datac";

dffeas \write_data_length[1] (
	.clk(altera_internal_jtag),
	.d(\header_in[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_data_length[0]~1_combout ),
	.q(\write_data_length[1]~q ),
	.prn(vcc));
defparam \write_data_length[1] .is_wysiwyg = "true";
defparam \write_data_length[1] .power_up = "low";

dffeas \write_data_length[2] (
	.clk(altera_internal_jtag),
	.d(altera_internal_jtag1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_data_length[0]~1_combout ),
	.q(\write_data_length[2]~q ),
	.prn(vcc));
defparam \write_data_length[2] .is_wysiwyg = "true";
defparam \write_data_length[2] .power_up = "low";

fiftyfivenm_lcell_comb \valid_write_data_length_byte_counter~11 (
	.dataa(\valid_write_data_length_byte_counter~10_combout ),
	.datab(\write_data_length[1]~q ),
	.datac(\write_data_length[2]~q ),
	.datad(\scan_length[0]~q ),
	.cin(gnd),
	.combout(\valid_write_data_length_byte_counter~11_combout ),
	.cout());
defparam \valid_write_data_length_byte_counter~11 .lut_mask = 16'hBEFF;
defparam \valid_write_data_length_byte_counter~11 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add4~16 (
	.dataa(\valid_write_data_length_byte_counter[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add4~15 ),
	.combout(\Add4~16_combout ),
	.cout(\Add4~17 ));
defparam \Add4~16 .lut_mask = 16'h5AAF;
defparam \Add4~16 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \valid_write_data_length_byte_counter~12 (
	.dataa(\valid_write_data_length_byte_counter[5]~1_combout ),
	.datab(\valid_write_data_length_byte_counter~11_combout ),
	.datac(\always2~0_combout ),
	.datad(\Add4~16_combout ),
	.cin(gnd),
	.combout(\valid_write_data_length_byte_counter~12_combout ),
	.cout());
defparam \valid_write_data_length_byte_counter~12 .lut_mask = 16'hFFFE;
defparam \valid_write_data_length_byte_counter~12 .sum_lutc_input = "datac";

dffeas \valid_write_data_length_byte_counter[8] (
	.clk(altera_internal_jtag),
	.d(\valid_write_data_length_byte_counter~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\valid_write_data_length_byte_counter[0]~2_combout ),
	.q(\valid_write_data_length_byte_counter[8]~q ),
	.prn(vcc));
defparam \valid_write_data_length_byte_counter[8] .is_wysiwyg = "true";
defparam \valid_write_data_length_byte_counter[8] .power_up = "low";

fiftyfivenm_lcell_comb \valid_write_data_length_byte_counter~13 (
	.dataa(\write_data_length[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\always2~0_combout ),
	.cin(gnd),
	.combout(\valid_write_data_length_byte_counter~13_combout ),
	.cout());
defparam \valid_write_data_length_byte_counter~13 .lut_mask = 16'hAAFF;
defparam \valid_write_data_length_byte_counter~13 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add2~0 (
	.dataa(\scan_length[1]~q ),
	.datab(\scan_length[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add2~0_combout ),
	.cout(\Add2~1 ));
defparam \Add2~0 .lut_mask = 16'h66EE;
defparam \Add2~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \valid_write_data_length_byte_counter~14 (
	.dataa(\valid_write_data_length_byte_counter~13_combout ),
	.datab(\Add2~0_combout ),
	.datac(\write_data_length[0]~q ),
	.datad(\write_data_length[2]~q ),
	.cin(gnd),
	.combout(\valid_write_data_length_byte_counter~14_combout ),
	.cout());
defparam \valid_write_data_length_byte_counter~14 .lut_mask = 16'hEFFE;
defparam \valid_write_data_length_byte_counter~14 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add4~18 (
	.dataa(\valid_write_data_length_byte_counter[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add4~17 ),
	.combout(\Add4~18_combout ),
	.cout(\Add4~19 ));
defparam \Add4~18 .lut_mask = 16'h5A5F;
defparam \Add4~18 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \valid_write_data_length_byte_counter~15 (
	.dataa(\valid_write_data_length_byte_counter[5]~1_combout ),
	.datab(\valid_write_data_length_byte_counter~14_combout ),
	.datac(\always2~0_combout ),
	.datad(\Add4~18_combout ),
	.cin(gnd),
	.combout(\valid_write_data_length_byte_counter~15_combout ),
	.cout());
defparam \valid_write_data_length_byte_counter~15 .lut_mask = 16'hFFFE;
defparam \valid_write_data_length_byte_counter~15 .sum_lutc_input = "datac";

dffeas \valid_write_data_length_byte_counter[9] (
	.clk(altera_internal_jtag),
	.d(\valid_write_data_length_byte_counter~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\valid_write_data_length_byte_counter[0]~2_combout ),
	.q(\valid_write_data_length_byte_counter[9]~q ),
	.prn(vcc));
defparam \valid_write_data_length_byte_counter[9] .is_wysiwyg = "true";
defparam \valid_write_data_length_byte_counter[9] .power_up = "low";

fiftyfivenm_lcell_comb \Add2~2 (
	.dataa(\scan_length[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~1 ),
	.combout(\Add2~2_combout ),
	.cout(\Add2~3 ));
defparam \Add2~2 .lut_mask = 16'h5A5F;
defparam \Add2~2 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \valid_write_data_length_byte_counter~16 (
	.dataa(\valid_write_data_length_byte_counter~10_combout ),
	.datab(\write_data_length[1]~q ),
	.datac(\Add2~2_combout ),
	.datad(\write_data_length[2]~q ),
	.cin(gnd),
	.combout(\valid_write_data_length_byte_counter~16_combout ),
	.cout());
defparam \valid_write_data_length_byte_counter~16 .lut_mask = 16'hFEFF;
defparam \valid_write_data_length_byte_counter~16 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add4~20 (
	.dataa(\valid_write_data_length_byte_counter[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add4~19 ),
	.combout(\Add4~20_combout ),
	.cout(\Add4~21 ));
defparam \Add4~20 .lut_mask = 16'h5AAF;
defparam \Add4~20 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \valid_write_data_length_byte_counter~17 (
	.dataa(\valid_write_data_length_byte_counter[5]~1_combout ),
	.datab(\valid_write_data_length_byte_counter~16_combout ),
	.datac(\always2~0_combout ),
	.datad(\Add4~20_combout ),
	.cin(gnd),
	.combout(\valid_write_data_length_byte_counter~17_combout ),
	.cout());
defparam \valid_write_data_length_byte_counter~17 .lut_mask = 16'hFFFE;
defparam \valid_write_data_length_byte_counter~17 .sum_lutc_input = "datac";

dffeas \valid_write_data_length_byte_counter[10] (
	.clk(altera_internal_jtag),
	.d(\valid_write_data_length_byte_counter~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\valid_write_data_length_byte_counter[0]~2_combout ),
	.q(\valid_write_data_length_byte_counter[10]~q ),
	.prn(vcc));
defparam \valid_write_data_length_byte_counter[10] .is_wysiwyg = "true";
defparam \valid_write_data_length_byte_counter[10] .power_up = "low";

fiftyfivenm_lcell_comb \Add4~22 (
	.dataa(\valid_write_data_length_byte_counter[11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add4~21 ),
	.combout(\Add4~22_combout ),
	.cout(\Add4~23 ));
defparam \Add4~22 .lut_mask = 16'h5A5F;
defparam \Add4~22 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add2~4 (
	.dataa(\scan_length[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~3 ),
	.combout(\Add2~4_combout ),
	.cout(\Add2~5 ));
defparam \Add2~4 .lut_mask = 16'h5AAF;
defparam \Add2~4 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \valid_write_data_length_byte_counter~18 (
	.dataa(\write_data_length[2]~q ),
	.datab(\Add2~4_combout ),
	.datac(\write_data_length[0]~q ),
	.datad(\write_data_length[1]~q ),
	.cin(gnd),
	.combout(\valid_write_data_length_byte_counter~18_combout ),
	.cout());
defparam \valid_write_data_length_byte_counter~18 .lut_mask = 16'hEFFE;
defparam \valid_write_data_length_byte_counter~18 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \valid_write_data_length_byte_counter~19 (
	.dataa(\valid_write_data_length_byte_counter[5]~1_combout ),
	.datab(\Add4~22_combout ),
	.datac(\always2~0_combout ),
	.datad(\valid_write_data_length_byte_counter~18_combout ),
	.cin(gnd),
	.combout(\valid_write_data_length_byte_counter~19_combout ),
	.cout());
defparam \valid_write_data_length_byte_counter~19 .lut_mask = 16'hFFAC;
defparam \valid_write_data_length_byte_counter~19 .sum_lutc_input = "datac";

dffeas \valid_write_data_length_byte_counter[11] (
	.clk(altera_internal_jtag),
	.d(\valid_write_data_length_byte_counter~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\valid_write_data_length_byte_counter[0]~2_combout ),
	.q(\valid_write_data_length_byte_counter[11]~q ),
	.prn(vcc));
defparam \valid_write_data_length_byte_counter[11] .is_wysiwyg = "true";
defparam \valid_write_data_length_byte_counter[11] .power_up = "low";

fiftyfivenm_lcell_comb \Equal13~2 (
	.dataa(\valid_write_data_length_byte_counter[8]~q ),
	.datab(\valid_write_data_length_byte_counter[9]~q ),
	.datac(\valid_write_data_length_byte_counter[10]~q ),
	.datad(\valid_write_data_length_byte_counter[11]~q ),
	.cin(gnd),
	.combout(\Equal13~2_combout ),
	.cout());
defparam \Equal13~2 .lut_mask = 16'h7FFF;
defparam \Equal13~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add2~6 (
	.dataa(\scan_length[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~5 ),
	.combout(\Add2~6_combout ),
	.cout(\Add2~7 ));
defparam \Add2~6 .lut_mask = 16'h5A5F;
defparam \Add2~6 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \valid_write_data_length_byte_counter~20 (
	.dataa(\valid_write_data_length_byte_counter~10_combout ),
	.datab(\write_data_length[2]~q ),
	.datac(\Add2~6_combout ),
	.datad(\write_data_length[1]~q ),
	.cin(gnd),
	.combout(\valid_write_data_length_byte_counter~20_combout ),
	.cout());
defparam \valid_write_data_length_byte_counter~20 .lut_mask = 16'hFEFF;
defparam \valid_write_data_length_byte_counter~20 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add4~24 (
	.dataa(\valid_write_data_length_byte_counter[12]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add4~23 ),
	.combout(\Add4~24_combout ),
	.cout(\Add4~25 ));
defparam \Add4~24 .lut_mask = 16'h5AAF;
defparam \Add4~24 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \valid_write_data_length_byte_counter~21 (
	.dataa(\valid_write_data_length_byte_counter[5]~1_combout ),
	.datab(\valid_write_data_length_byte_counter~20_combout ),
	.datac(\always2~0_combout ),
	.datad(\Add4~24_combout ),
	.cin(gnd),
	.combout(\valid_write_data_length_byte_counter~21_combout ),
	.cout());
defparam \valid_write_data_length_byte_counter~21 .lut_mask = 16'hFFFE;
defparam \valid_write_data_length_byte_counter~21 .sum_lutc_input = "datac";

dffeas \valid_write_data_length_byte_counter[12] (
	.clk(altera_internal_jtag),
	.d(\valid_write_data_length_byte_counter~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\valid_write_data_length_byte_counter[0]~2_combout ),
	.q(\valid_write_data_length_byte_counter[12]~q ),
	.prn(vcc));
defparam \valid_write_data_length_byte_counter[12] .is_wysiwyg = "true";
defparam \valid_write_data_length_byte_counter[12] .power_up = "low";

fiftyfivenm_lcell_comb \Add2~8 (
	.dataa(\scan_length[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~7 ),
	.combout(\Add2~8_combout ),
	.cout(\Add2~9 ));
defparam \Add2~8 .lut_mask = 16'h5AAF;
defparam \Add2~8 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \valid_write_data_length_byte_counter~22 (
	.dataa(\write_data_length[2]~q ),
	.datab(\valid_write_data_length_byte_counter~13_combout ),
	.datac(\Add2~8_combout ),
	.datad(\write_data_length[0]~q ),
	.cin(gnd),
	.combout(\valid_write_data_length_byte_counter~22_combout ),
	.cout());
defparam \valid_write_data_length_byte_counter~22 .lut_mask = 16'hFEFF;
defparam \valid_write_data_length_byte_counter~22 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add4~26 (
	.dataa(\valid_write_data_length_byte_counter[13]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add4~25 ),
	.combout(\Add4~26_combout ),
	.cout(\Add4~27 ));
defparam \Add4~26 .lut_mask = 16'h5A5F;
defparam \Add4~26 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \valid_write_data_length_byte_counter~23 (
	.dataa(\valid_write_data_length_byte_counter[5]~1_combout ),
	.datab(\valid_write_data_length_byte_counter~22_combout ),
	.datac(\always2~0_combout ),
	.datad(\Add4~26_combout ),
	.cin(gnd),
	.combout(\valid_write_data_length_byte_counter~23_combout ),
	.cout());
defparam \valid_write_data_length_byte_counter~23 .lut_mask = 16'hFFFE;
defparam \valid_write_data_length_byte_counter~23 .sum_lutc_input = "datac";

dffeas \valid_write_data_length_byte_counter[13] (
	.clk(altera_internal_jtag),
	.d(\valid_write_data_length_byte_counter~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\valid_write_data_length_byte_counter[0]~2_combout ),
	.q(\valid_write_data_length_byte_counter[13]~q ),
	.prn(vcc));
defparam \valid_write_data_length_byte_counter[13] .is_wysiwyg = "true";
defparam \valid_write_data_length_byte_counter[13] .power_up = "low";

fiftyfivenm_lcell_comb \Add2~10 (
	.dataa(\scan_length[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~9 ),
	.combout(\Add2~10_combout ),
	.cout(\Add2~11 ));
defparam \Add2~10 .lut_mask = 16'h5A5F;
defparam \Add2~10 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \valid_write_data_length_byte_counter~24 (
	.dataa(\write_data_length[0]~q ),
	.datab(\write_data_length[1]~q ),
	.datac(\write_data_length[2]~q ),
	.datad(\always2~0_combout ),
	.cin(gnd),
	.combout(\valid_write_data_length_byte_counter~24_combout ),
	.cout());
defparam \valid_write_data_length_byte_counter~24 .lut_mask = 16'hFEFF;
defparam \valid_write_data_length_byte_counter~24 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \valid_write_data_length_byte_counter~25 (
	.dataa(\Add2~10_combout ),
	.datab(\valid_write_data_length_byte_counter~24_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\valid_write_data_length_byte_counter~25_combout ),
	.cout());
defparam \valid_write_data_length_byte_counter~25 .lut_mask = 16'hEEEE;
defparam \valid_write_data_length_byte_counter~25 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add4~28 (
	.dataa(\valid_write_data_length_byte_counter[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add4~27 ),
	.combout(\Add4~28_combout ),
	.cout(\Add4~29 ));
defparam \Add4~28 .lut_mask = 16'h5AAF;
defparam \Add4~28 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \valid_write_data_length_byte_counter~26 (
	.dataa(\valid_write_data_length_byte_counter[5]~1_combout ),
	.datab(\valid_write_data_length_byte_counter~25_combout ),
	.datac(\always2~0_combout ),
	.datad(\Add4~28_combout ),
	.cin(gnd),
	.combout(\valid_write_data_length_byte_counter~26_combout ),
	.cout());
defparam \valid_write_data_length_byte_counter~26 .lut_mask = 16'hFFFE;
defparam \valid_write_data_length_byte_counter~26 .sum_lutc_input = "datac";

dffeas \valid_write_data_length_byte_counter[14] (
	.clk(altera_internal_jtag),
	.d(\valid_write_data_length_byte_counter~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\valid_write_data_length_byte_counter[0]~2_combout ),
	.q(\valid_write_data_length_byte_counter[14]~q ),
	.prn(vcc));
defparam \valid_write_data_length_byte_counter[14] .is_wysiwyg = "true";
defparam \valid_write_data_length_byte_counter[14] .power_up = "low";

fiftyfivenm_lcell_comb \Add4~30 (
	.dataa(\valid_write_data_length_byte_counter[15]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add4~29 ),
	.combout(\Add4~30_combout ),
	.cout(\Add4~31 ));
defparam \Add4~30 .lut_mask = 16'h5A5F;
defparam \Add4~30 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add2~12 (
	.dataa(\scan_length[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~11 ),
	.combout(\Add2~12_combout ),
	.cout(\Add2~13 ));
defparam \Add2~12 .lut_mask = 16'h5AAF;
defparam \Add2~12 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \valid_write_data_length_byte_counter~27 (
	.dataa(\Add2~12_combout ),
	.datab(\valid_write_data_length_byte_counter~24_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\valid_write_data_length_byte_counter~27_combout ),
	.cout());
defparam \valid_write_data_length_byte_counter~27 .lut_mask = 16'hEEEE;
defparam \valid_write_data_length_byte_counter~27 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \valid_write_data_length_byte_counter~28 (
	.dataa(\valid_write_data_length_byte_counter[5]~1_combout ),
	.datab(\always2~0_combout ),
	.datac(\Add4~30_combout ),
	.datad(\valid_write_data_length_byte_counter~27_combout ),
	.cin(gnd),
	.combout(\valid_write_data_length_byte_counter~28_combout ),
	.cout());
defparam \valid_write_data_length_byte_counter~28 .lut_mask = 16'hFFFE;
defparam \valid_write_data_length_byte_counter~28 .sum_lutc_input = "datac";

dffeas \valid_write_data_length_byte_counter[15] (
	.clk(altera_internal_jtag),
	.d(\valid_write_data_length_byte_counter~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\valid_write_data_length_byte_counter[0]~2_combout ),
	.q(\valid_write_data_length_byte_counter[15]~q ),
	.prn(vcc));
defparam \valid_write_data_length_byte_counter[15] .is_wysiwyg = "true";
defparam \valid_write_data_length_byte_counter[15] .power_up = "low";

fiftyfivenm_lcell_comb \Equal13~3 (
	.dataa(\valid_write_data_length_byte_counter[12]~q ),
	.datab(\valid_write_data_length_byte_counter[13]~q ),
	.datac(\valid_write_data_length_byte_counter[14]~q ),
	.datad(\valid_write_data_length_byte_counter[15]~q ),
	.cin(gnd),
	.combout(\Equal13~3_combout ),
	.cout());
defparam \Equal13~3 .lut_mask = 16'h7FFF;
defparam \Equal13~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Equal13~4 (
	.dataa(\Equal13~0_combout ),
	.datab(\Equal13~1_combout ),
	.datac(\Equal13~2_combout ),
	.datad(\Equal13~3_combout ),
	.cin(gnd),
	.combout(\Equal13~4_combout ),
	.cout());
defparam \Equal13~4 .lut_mask = 16'hFFFE;
defparam \Equal13~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add4~32 (
	.dataa(\valid_write_data_length_byte_counter[16]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add4~31 ),
	.combout(\Add4~32_combout ),
	.cout(\Add4~33 ));
defparam \Add4~32 .lut_mask = 16'h5AAF;
defparam \Add4~32 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add2~14 (
	.dataa(\scan_length[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~13 ),
	.combout(\Add2~14_combout ),
	.cout(\Add2~15 ));
defparam \Add2~14 .lut_mask = 16'h5A5F;
defparam \Add2~14 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \valid_write_data_length_byte_counter~29 (
	.dataa(\Add2~14_combout ),
	.datab(\valid_write_data_length_byte_counter~24_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\valid_write_data_length_byte_counter~29_combout ),
	.cout());
defparam \valid_write_data_length_byte_counter~29 .lut_mask = 16'hEEEE;
defparam \valid_write_data_length_byte_counter~29 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \valid_write_data_length_byte_counter~30 (
	.dataa(\valid_write_data_length_byte_counter[5]~1_combout ),
	.datab(\always2~0_combout ),
	.datac(\Add4~32_combout ),
	.datad(\valid_write_data_length_byte_counter~29_combout ),
	.cin(gnd),
	.combout(\valid_write_data_length_byte_counter~30_combout ),
	.cout());
defparam \valid_write_data_length_byte_counter~30 .lut_mask = 16'hFFFE;
defparam \valid_write_data_length_byte_counter~30 .sum_lutc_input = "datac";

dffeas \valid_write_data_length_byte_counter[16] (
	.clk(altera_internal_jtag),
	.d(\valid_write_data_length_byte_counter~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\valid_write_data_length_byte_counter[0]~2_combout ),
	.q(\valid_write_data_length_byte_counter[16]~q ),
	.prn(vcc));
defparam \valid_write_data_length_byte_counter[16] .is_wysiwyg = "true";
defparam \valid_write_data_length_byte_counter[16] .power_up = "low";

fiftyfivenm_lcell_comb \Add4~34 (
	.dataa(\valid_write_data_length_byte_counter[17]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add4~33 ),
	.combout(\Add4~34_combout ),
	.cout(\Add4~35 ));
defparam \Add4~34 .lut_mask = 16'h5A5F;
defparam \Add4~34 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \Add2~16 (
	.dataa(\scan_length[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~15 ),
	.combout(\Add2~16_combout ),
	.cout(\Add2~17 ));
defparam \Add2~16 .lut_mask = 16'h5AAF;
defparam \Add2~16 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \valid_write_data_length_byte_counter~31 (
	.dataa(\valid_write_data_length_byte_counter~24_combout ),
	.datab(\Add2~16_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\valid_write_data_length_byte_counter~31_combout ),
	.cout());
defparam \valid_write_data_length_byte_counter~31 .lut_mask = 16'hEEEE;
defparam \valid_write_data_length_byte_counter~31 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \valid_write_data_length_byte_counter~32 (
	.dataa(\valid_write_data_length_byte_counter[5]~1_combout ),
	.datab(\always2~0_combout ),
	.datac(\Add4~34_combout ),
	.datad(\valid_write_data_length_byte_counter~31_combout ),
	.cin(gnd),
	.combout(\valid_write_data_length_byte_counter~32_combout ),
	.cout());
defparam \valid_write_data_length_byte_counter~32 .lut_mask = 16'hFFFE;
defparam \valid_write_data_length_byte_counter~32 .sum_lutc_input = "datac";

dffeas \valid_write_data_length_byte_counter[17] (
	.clk(altera_internal_jtag),
	.d(\valid_write_data_length_byte_counter~32_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\valid_write_data_length_byte_counter[0]~2_combout ),
	.q(\valid_write_data_length_byte_counter[17]~q ),
	.prn(vcc));
defparam \valid_write_data_length_byte_counter[17] .is_wysiwyg = "true";
defparam \valid_write_data_length_byte_counter[17] .power_up = "low";

fiftyfivenm_lcell_comb \Add2~18 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add2~17 ),
	.combout(\Add2~18_combout ),
	.cout());
defparam \Add2~18 .lut_mask = 16'hF0F0;
defparam \Add2~18 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \valid_write_data_length_byte_counter~33 (
	.dataa(\valid_write_data_length_byte_counter~24_combout ),
	.datab(\Add2~18_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\valid_write_data_length_byte_counter~33_combout ),
	.cout());
defparam \valid_write_data_length_byte_counter~33 .lut_mask = 16'hEEEE;
defparam \valid_write_data_length_byte_counter~33 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Add4~36 (
	.dataa(\valid_write_data_length_byte_counter[18]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add4~35 ),
	.combout(\Add4~36_combout ),
	.cout());
defparam \Add4~36 .lut_mask = 16'h5A5A;
defparam \Add4~36 .sum_lutc_input = "cin";

fiftyfivenm_lcell_comb \valid_write_data_length_byte_counter~34 (
	.dataa(\valid_write_data_length_byte_counter[5]~1_combout ),
	.datab(\valid_write_data_length_byte_counter~33_combout ),
	.datac(\always2~0_combout ),
	.datad(\Add4~36_combout ),
	.cin(gnd),
	.combout(\valid_write_data_length_byte_counter~34_combout ),
	.cout());
defparam \valid_write_data_length_byte_counter~34 .lut_mask = 16'hFFFE;
defparam \valid_write_data_length_byte_counter~34 .sum_lutc_input = "datac";

dffeas \valid_write_data_length_byte_counter[18] (
	.clk(altera_internal_jtag),
	.d(\valid_write_data_length_byte_counter~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\valid_write_data_length_byte_counter[0]~2_combout ),
	.q(\valid_write_data_length_byte_counter[18]~q ),
	.prn(vcc));
defparam \valid_write_data_length_byte_counter[18] .is_wysiwyg = "true";
defparam \valid_write_data_length_byte_counter[18] .power_up = "low";

fiftyfivenm_lcell_comb \Equal13~5 (
	.dataa(\Equal13~4_combout ),
	.datab(\valid_write_data_length_byte_counter[16]~q ),
	.datac(\valid_write_data_length_byte_counter[17]~q ),
	.datad(\valid_write_data_length_byte_counter[18]~q ),
	.cin(gnd),
	.combout(\Equal13~5_combout ),
	.cout());
defparam \Equal13~5 .lut_mask = 16'hFFFD;
defparam \Equal13~5 .sum_lutc_input = "datac";

dffeas write_data_valid(
	.clk(altera_internal_jtag),
	.d(\Equal13~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dr_data_in[1]~0_combout ),
	.q(\write_data_valid~q ),
	.prn(vcc));
defparam write_data_valid.is_wysiwyg = "true";
defparam write_data_valid.power_up = "low";

fiftyfivenm_lcell_comb \write_data_bit_counter~0 (
	.dataa(\write_data_bit_counter[0]~q ),
	.datab(gnd),
	.datac(virtual_state_sdr),
	.datad(\write_state.ST_WRITE_DATA~q ),
	.cin(gnd),
	.combout(\write_data_bit_counter~0_combout ),
	.cout());
defparam \write_data_bit_counter~0 .lut_mask = 16'hFF5F;
defparam \write_data_bit_counter~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \write_data_bit_counter[0]~1 (
	.dataa(\Equal14~0_combout ),
	.datab(virtual_state_sdr),
	.datac(\write_state.ST_WRITE_DATA~q ),
	.datad(virtual_state_cdr),
	.cin(gnd),
	.combout(\write_data_bit_counter[0]~1_combout ),
	.cout());
defparam \write_data_bit_counter[0]~1 .lut_mask = 16'hFBFF;
defparam \write_data_bit_counter[0]~1 .sum_lutc_input = "datac";

dffeas \write_data_bit_counter[0] (
	.clk(altera_internal_jtag),
	.d(\write_data_bit_counter~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_data_bit_counter[0]~1_combout ),
	.q(\write_data_bit_counter[0]~q ),
	.prn(vcc));
defparam \write_data_bit_counter[0] .is_wysiwyg = "true";
defparam \write_data_bit_counter[0] .power_up = "low";

fiftyfivenm_lcell_comb \write_data_bit_counter~2 (
	.dataa(\write_data_bit_counter[0]~q ),
	.datab(\write_data_bit_counter[1]~q ),
	.datac(virtual_state_sdr),
	.datad(\write_state.ST_WRITE_DATA~q ),
	.cin(gnd),
	.combout(\write_data_bit_counter~2_combout ),
	.cout());
defparam \write_data_bit_counter~2 .lut_mask = 16'hFF6F;
defparam \write_data_bit_counter~2 .sum_lutc_input = "datac";

dffeas \write_data_bit_counter[1] (
	.clk(altera_internal_jtag),
	.d(\write_data_bit_counter~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_data_bit_counter[0]~1_combout ),
	.q(\write_data_bit_counter[1]~q ),
	.prn(vcc));
defparam \write_data_bit_counter[1] .is_wysiwyg = "true";
defparam \write_data_bit_counter[1] .power_up = "low";

fiftyfivenm_lcell_comb \Add3~0 (
	.dataa(gnd),
	.datab(\write_data_bit_counter[0]~q ),
	.datac(\write_data_bit_counter[1]~q ),
	.datad(\write_data_bit_counter[2]~q ),
	.cin(gnd),
	.combout(\Add3~0_combout ),
	.cout());
defparam \Add3~0 .lut_mask = 16'hC33C;
defparam \Add3~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \write_data_bit_counter~3 (
	.dataa(\Add3~0_combout ),
	.datab(gnd),
	.datac(virtual_state_sdr),
	.datad(\write_state.ST_WRITE_DATA~q ),
	.cin(gnd),
	.combout(\write_data_bit_counter~3_combout ),
	.cout());
defparam \write_data_bit_counter~3 .lut_mask = 16'hFF5F;
defparam \write_data_bit_counter~3 .sum_lutc_input = "datac";

dffeas \write_data_bit_counter[2] (
	.clk(altera_internal_jtag),
	.d(\write_data_bit_counter~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\write_data_bit_counter[0]~1_combout ),
	.q(\write_data_bit_counter[2]~q ),
	.prn(vcc));
defparam \write_data_bit_counter[2] .is_wysiwyg = "true";
defparam \write_data_bit_counter[2] .power_up = "low";

fiftyfivenm_lcell_comb \always2~0 (
	.dataa(\write_data_valid~q ),
	.datab(\write_data_bit_counter[0]~q ),
	.datac(\write_data_bit_counter[1]~q ),
	.datad(\write_data_bit_counter[2]~q ),
	.cin(gnd),
	.combout(\always2~0_combout ),
	.cout());
defparam \always2~0 .lut_mask = 16'hEFFF;
defparam \always2~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \idle_remover_sink_data[0]~0 (
	.dataa(virtual_state_sdr),
	.datab(\Equal14~0_combout ),
	.datac(\write_state.ST_WRITE_DATA~q ),
	.datad(\always2~0_combout ),
	.cin(gnd),
	.combout(\idle_remover_sink_data[0]~0_combout ),
	.cout());
defparam \idle_remover_sink_data[0]~0 .lut_mask = 16'hFFFD;
defparam \idle_remover_sink_data[0]~0 .sum_lutc_input = "datac";

dffeas \dr_data_in[3] (
	.clk(altera_internal_jtag),
	.d(\dr_data_in[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dr_data_in[1]~0_combout ),
	.q(\dr_data_in[3]~q ),
	.prn(vcc));
defparam \dr_data_in[3] .is_wysiwyg = "true";
defparam \dr_data_in[3] .power_up = "low";

dffeas \dr_data_in[2] (
	.clk(altera_internal_jtag),
	.d(\dr_data_in[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dr_data_in[1]~0_combout ),
	.q(\dr_data_in[2]~q ),
	.prn(vcc));
defparam \dr_data_in[2] .is_wysiwyg = "true";
defparam \dr_data_in[2] .power_up = "low";

dffeas \dr_data_in[1] (
	.clk(altera_internal_jtag),
	.d(\dr_data_in[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\dr_data_in[1]~0_combout ),
	.q(\dr_data_in[1]~q ),
	.prn(vcc));
defparam \dr_data_in[1] .is_wysiwyg = "true";
defparam \dr_data_in[1] .power_up = "low";

endmodule

module ADC_altera_avalon_st_idle_inserter (
	data1_0,
	data1_2,
	data1_1,
	data1_6,
	data1_7,
	data1_5,
	data1_3,
	data1_4,
	out_data,
	out_data1,
	full1,
	reset_n,
	idle_inserter_source_ready,
	in_ready,
	out_data2,
	clk)/* synthesis synthesis_greybox=1 */;
input 	data1_0;
input 	data1_2;
input 	data1_1;
input 	data1_6;
input 	data1_7;
input 	data1_5;
input 	data1_3;
input 	data1_4;
output 	out_data;
output 	out_data1;
input 	full1;
input 	reset_n;
input 	idle_inserter_source_ready;
output 	in_ready;
output 	out_data2;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \out_data~0_combout ;
wire \received_esc~0_combout ;
wire \received_esc~q ;
wire \out_data~1_combout ;


fiftyfivenm_lcell_comb \out_data~2 (
	.dataa(\out_data~0_combout ),
	.datab(\out_data~1_combout ),
	.datac(data1_3),
	.datad(data1_4),
	.cin(gnd),
	.combout(out_data),
	.cout());
defparam \out_data~2 .lut_mask = 16'hFEFF;
defparam \out_data~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data~3 (
	.dataa(data1_0),
	.datab(out_data),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_data1),
	.cout());
defparam \out_data~3 .lut_mask = 16'hEEEE;
defparam \out_data~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \in_ready~0 (
	.dataa(idle_inserter_source_ready),
	.datab(gnd),
	.datac(out_data),
	.datad(full1),
	.cin(gnd),
	.combout(in_ready),
	.cout());
defparam \in_ready~0 .lut_mask = 16'hAFFF;
defparam \in_ready~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\received_esc~q ),
	.datad(data1_5),
	.cin(gnd),
	.combout(out_data2),
	.cout());
defparam \out_data~4 .lut_mask = 16'h0FF0;
defparam \out_data~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data~0 (
	.dataa(gnd),
	.datab(data1_0),
	.datac(data1_2),
	.datad(data1_1),
	.cin(gnd),
	.combout(\out_data~0_combout ),
	.cout());
defparam \out_data~0 .lut_mask = 16'hC33C;
defparam \out_data~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \received_esc~0 (
	.dataa(out_data),
	.datab(\received_esc~q ),
	.datac(full1),
	.datad(idle_inserter_source_ready),
	.cin(gnd),
	.combout(\received_esc~0_combout ),
	.cout());
defparam \received_esc~0 .lut_mask = 16'hEFFE;
defparam \received_esc~0 .sum_lutc_input = "datac";

dffeas received_esc(
	.clk(clk),
	.d(\received_esc~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\received_esc~q ),
	.prn(vcc));
defparam received_esc.is_wysiwyg = "true";
defparam received_esc.power_up = "low";

fiftyfivenm_lcell_comb \out_data~1 (
	.dataa(data1_6),
	.datab(\received_esc~q ),
	.datac(data1_7),
	.datad(data1_5),
	.cin(gnd),
	.combout(\out_data~1_combout ),
	.cout());
defparam \out_data~1 .lut_mask = 16'hBFFF;
defparam \out_data~1 .sum_lutc_input = "datac";

endmodule

module ADC_altera_avalon_st_idle_remover (
	reset_n,
	idle_remover_sink_data_3,
	idle_remover_sink_valid,
	idle_remover_sink_data_7,
	idle_remover_sink_data_6,
	idle_remover_sink_data_4,
	idle_remover_sink_data_5,
	idle_remover_sink_data_1,
	idle_remover_sink_data_0,
	idle_remover_sink_data_2,
	out_data_5,
	out_valid1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset_n;
input 	idle_remover_sink_data_3;
input 	idle_remover_sink_valid;
input 	idle_remover_sink_data_7;
input 	idle_remover_sink_data_6;
input 	idle_remover_sink_data_4;
input 	idle_remover_sink_data_5;
input 	idle_remover_sink_data_1;
input 	idle_remover_sink_data_0;
input 	idle_remover_sink_data_2;
output 	out_data_5;
output 	out_valid1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \out_valid~3_combout ;
wire \Equal0~0_combout ;
wire \out_valid~4_combout ;
wire \Equal0~1_combout ;
wire \out_valid~2_combout ;
wire \received_esc~0_combout ;
wire \received_esc~q ;


fiftyfivenm_lcell_comb \out_data[5]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(idle_remover_sink_data_5),
	.datad(\received_esc~q ),
	.cin(gnd),
	.combout(out_data_5),
	.cout());
defparam \out_data[5]~0 .lut_mask = 16'h0FF0;
defparam \out_data[5]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb out_valid(
	.dataa(idle_remover_sink_data_7),
	.datab(\out_valid~3_combout ),
	.datac(\Equal0~0_combout ),
	.datad(\out_valid~2_combout ),
	.cin(gnd),
	.combout(out_valid1),
	.cout());
defparam out_valid.lut_mask = 16'hFFEF;
defparam out_valid.sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_valid~3 (
	.dataa(idle_remover_sink_data_1),
	.datab(\received_esc~q ),
	.datac(idle_remover_sink_data_0),
	.datad(idle_remover_sink_data_2),
	.cin(gnd),
	.combout(\out_valid~3_combout ),
	.cout());
defparam \out_valid~3 .lut_mask = 16'hEFFF;
defparam \out_valid~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Equal0~0 (
	.dataa(idle_remover_sink_data_3),
	.datab(idle_remover_sink_data_6),
	.datac(idle_remover_sink_data_4),
	.datad(idle_remover_sink_data_5),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'hEFFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_valid~4 (
	.dataa(idle_remover_sink_data_7),
	.datab(\out_valid~3_combout ),
	.datac(gnd),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\out_valid~4_combout ),
	.cout());
defparam \out_valid~4 .lut_mask = 16'hEEFF;
defparam \out_valid~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Equal0~1 (
	.dataa(idle_remover_sink_data_1),
	.datab(gnd),
	.datac(idle_remover_sink_data_0),
	.datad(idle_remover_sink_data_2),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'hAFFF;
defparam \Equal0~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_valid~2 (
	.dataa(idle_remover_sink_valid),
	.datab(idle_remover_sink_data_7),
	.datac(\Equal0~0_combout ),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(\out_valid~2_combout ),
	.cout());
defparam \out_valid~2 .lut_mask = 16'hEFFF;
defparam \out_valid~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \received_esc~0 (
	.dataa(idle_remover_sink_valid),
	.datab(\received_esc~q ),
	.datac(\out_valid~4_combout ),
	.datad(\out_valid~2_combout ),
	.cin(gnd),
	.combout(\received_esc~0_combout ),
	.cout());
defparam \received_esc~0 .lut_mask = 16'hEFFF;
defparam \received_esc~0 .sum_lutc_input = "datac";

dffeas received_esc(
	.clk(clk),
	.d(\received_esc~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\received_esc~q ),
	.prn(vcc));
defparam received_esc.is_wysiwyg = "true";
defparam received_esc.power_up = "low";

endmodule

module ADC_altera_std_synchronizer_3 (
	dreg_6,
	reset_n,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_6;
input 	reset_n;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;
wire \dreg[1]~q ;
wire \dreg[2]~q ;
wire \dreg[3]~q ;
wire \dreg[4]~q ;
wire \dreg[5]~q ;


dffeas \dreg[6] (
	.clk(clk),
	.d(\dreg[5]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_6),
	.prn(vcc));
defparam \dreg[6] .is_wysiwyg = "true";
defparam \dreg[6] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[1]~q ),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas \dreg[2] (
	.clk(clk),
	.d(\dreg[1]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[2]~q ),
	.prn(vcc));
defparam \dreg[2] .is_wysiwyg = "true";
defparam \dreg[2] .power_up = "low";

dffeas \dreg[3] (
	.clk(clk),
	.d(\dreg[2]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[3]~q ),
	.prn(vcc));
defparam \dreg[3] .is_wysiwyg = "true";
defparam \dreg[3] .power_up = "low";

dffeas \dreg[4] (
	.clk(clk),
	.d(\dreg[3]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[4]~q ),
	.prn(vcc));
defparam \dreg[4] .is_wysiwyg = "true";
defparam \dreg[4] .power_up = "low";

dffeas \dreg[5] (
	.clk(clk),
	.d(\dreg[4]~q ),
	.asdata(vcc),
	.clrn(!reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[5]~q ),
	.prn(vcc));
defparam \dreg[5] .is_wysiwyg = "true";
defparam \dreg[5] .power_up = "low";

endmodule

module ADC_altera_std_synchronizer_4 (
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module ADC_altera_std_synchronizer_5 (
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module ADC_altera_std_synchronizer_6 (
	dreg_1,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module ADC_altera_std_synchronizer_7 (
	dreg_1,
	reset_n,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_1;
input 	reset_n;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;
wire \dreg[0]~q ;


dffeas \dreg[1] (
	.clk(clk),
	.d(\dreg[0]~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_1),
	.prn(vcc));
defparam \dreg[1] .is_wysiwyg = "true";
defparam \dreg[1] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\dreg[0]~q ),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

endmodule

module ADC_altera_jtag_sld_node (
	virtual_state_sdr,
	virtual_state_cdr,
	virtual_state_udr,
	state_4,
	splitter_nodes_receive_0_3,
	virtual_ir_scan_reg,
	state_3,
	state_8)/* synthesis synthesis_greybox=1 */;
output 	virtual_state_sdr;
output 	virtual_state_cdr;
output 	virtual_state_udr;
input 	state_4;
input 	splitter_nodes_receive_0_3;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ADC_sld_virtual_jtag_basic_1 sld_virtual_jtag_component(
	.virtual_state_sdr(virtual_state_sdr),
	.virtual_state_cdr1(virtual_state_cdr),
	.virtual_state_udr1(virtual_state_udr),
	.state_4(state_4),
	.splitter_nodes_receive_0_3(splitter_nodes_receive_0_3),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8));

endmodule

module ADC_sld_virtual_jtag_basic_1 (
	virtual_state_sdr,
	virtual_state_cdr1,
	virtual_state_udr1,
	state_4,
	splitter_nodes_receive_0_3,
	virtual_ir_scan_reg,
	state_3,
	state_8)/* synthesis synthesis_greybox=1 */;
output 	virtual_state_sdr;
output 	virtual_state_cdr1;
output 	virtual_state_udr1;
input 	state_4;
input 	splitter_nodes_receive_0_3;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fiftyfivenm_lcell_comb \virtual_state_sdr~0 (
	.dataa(splitter_nodes_receive_0_3),
	.datab(state_4),
	.datac(gnd),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(virtual_state_sdr),
	.cout());
defparam \virtual_state_sdr~0 .lut_mask = 16'hFF77;
defparam \virtual_state_sdr~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb virtual_state_cdr(
	.dataa(virtual_ir_scan_reg),
	.datab(gnd),
	.datac(splitter_nodes_receive_0_3),
	.datad(state_3),
	.cin(gnd),
	.combout(virtual_state_cdr1),
	.cout());
defparam virtual_state_cdr.lut_mask = 16'hAFFF;
defparam virtual_state_cdr.sum_lutc_input = "datac";

fiftyfivenm_lcell_comb virtual_state_udr(
	.dataa(splitter_nodes_receive_0_3),
	.datab(state_8),
	.datac(gnd),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(virtual_state_udr1),
	.cout());
defparam virtual_state_udr.lut_mask = 16'hEEFF;
defparam virtual_state_udr.sum_lutc_input = "datac";

endmodule

module ADC_altera_avalon_st_packets_to_bytes (
	out_endofpacket,
	reset_n,
	out_data_0,
	out_valid1,
	in_data_toggle,
	dreg_6,
	out_data_2,
	out_data_1,
	out_data_6,
	out_data_7,
	out_data_5,
	out_data_3,
	out_data_4,
	out_data_01,
	out_startofpacket,
	out_data_21,
	out_data_11,
	out_data_51,
	out_data_71,
	out_data_61,
	out_data_41,
	out_data_31,
	out_valid2,
	in_ready1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	out_endofpacket;
input 	reset_n;
output 	out_data_0;
output 	out_valid1;
input 	in_data_toggle;
input 	dreg_6;
output 	out_data_2;
output 	out_data_1;
output 	out_data_6;
output 	out_data_7;
output 	out_data_5;
output 	out_data_3;
output 	out_data_4;
input 	out_data_01;
input 	out_startofpacket;
input 	out_data_21;
input 	out_data_11;
input 	out_data_51;
input 	out_data_71;
input 	out_data_61;
input 	out_data_41;
input 	out_data_31;
input 	out_valid2;
output 	in_ready1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \in_ready~2_combout ;
wire \sent_esc~0_combout ;
wire \sent_esc~q ;
wire \in_ready~0_combout ;
wire \in_ready~1_combout ;
wire \in_ready~3_combout ;
wire \sent_channel_char~0_combout ;
wire \sent_channel_char~q ;
wire \sent_channel~0_combout ;
wire \sent_channel~1_combout ;
wire \sent_channel~q ;
wire \stored_channel[0]~0_combout ;
wire \stored_channel[0]~q ;
wire \always0~0_combout ;
wire \in_ready~4_combout ;
wire \sent_eop~2_combout ;
wire \sent_eop~q ;
wire \always0~2_combout ;
wire \sent_sop~3_combout ;
wire \sent_sop~2_combout ;
wire \sent_sop~q ;
wire \out_data[7]~0_combout ;
wire \out_data[7]~1_combout ;
wire \always0~1_combout ;
wire \out_data~2_combout ;
wire \out_valid~0_combout ;
wire \out_data~3_combout ;
wire \out_data~4_combout ;
wire \out_data~5_combout ;
wire \out_data~6_combout ;
wire \out_data~7_combout ;
wire \out_data~8_combout ;
wire \out_data~9_combout ;
wire \out_data~10_combout ;
wire \out_data~11_combout ;


dffeas \out_data[0] (
	.clk(clk),
	.d(\out_data~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~2_combout ),
	.q(out_data_0),
	.prn(vcc));
defparam \out_data[0] .is_wysiwyg = "true";
defparam \out_data[0] .power_up = "low";

dffeas out_valid(
	.clk(clk),
	.d(\out_valid~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_valid1),
	.prn(vcc));
defparam out_valid.is_wysiwyg = "true";
defparam out_valid.power_up = "low";

dffeas \out_data[2] (
	.clk(clk),
	.d(\out_data~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~2_combout ),
	.q(out_data_2),
	.prn(vcc));
defparam \out_data[2] .is_wysiwyg = "true";
defparam \out_data[2] .power_up = "low";

dffeas \out_data[1] (
	.clk(clk),
	.d(\out_data~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~2_combout ),
	.q(out_data_1),
	.prn(vcc));
defparam \out_data[1] .is_wysiwyg = "true";
defparam \out_data[1] .power_up = "low";

dffeas \out_data[6] (
	.clk(clk),
	.d(\out_data~6_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~2_combout ),
	.q(out_data_6),
	.prn(vcc));
defparam \out_data[6] .is_wysiwyg = "true";
defparam \out_data[6] .power_up = "low";

dffeas \out_data[7] (
	.clk(clk),
	.d(\out_data~7_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~2_combout ),
	.q(out_data_7),
	.prn(vcc));
defparam \out_data[7] .is_wysiwyg = "true";
defparam \out_data[7] .power_up = "low";

dffeas \out_data[5] (
	.clk(clk),
	.d(\out_data~9_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~2_combout ),
	.q(out_data_5),
	.prn(vcc));
defparam \out_data[5] .is_wysiwyg = "true";
defparam \out_data[5] .power_up = "low";

dffeas \out_data[3] (
	.clk(clk),
	.d(\out_data~10_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~2_combout ),
	.q(out_data_3),
	.prn(vcc));
defparam \out_data[3] .is_wysiwyg = "true";
defparam \out_data[3] .power_up = "low";

dffeas \out_data[4] (
	.clk(clk),
	.d(\out_data~11_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~2_combout ),
	.q(out_data_4),
	.prn(vcc));
defparam \out_data[4] .is_wysiwyg = "true";
defparam \out_data[4] .power_up = "low";

fiftyfivenm_lcell_comb in_ready(
	.dataa(\in_ready~4_combout ),
	.datab(\in_ready~0_combout ),
	.datac(\in_ready~1_combout ),
	.datad(\always0~2_combout ),
	.cin(gnd),
	.combout(in_ready1),
	.cout());
defparam in_ready.lut_mask = 16'hFEFF;
defparam in_ready.sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \in_ready~2 (
	.dataa(out_valid2),
	.datab(in_data_toggle),
	.datac(dreg_6),
	.datad(out_valid1),
	.cin(gnd),
	.combout(\in_ready~2_combout ),
	.cout());
defparam \in_ready~2 .lut_mask = 16'hBEFF;
defparam \in_ready~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \sent_esc~0 (
	.dataa(\sent_esc~q ),
	.datab(\always0~2_combout ),
	.datac(\in_ready~4_combout ),
	.datad(\in_ready~3_combout ),
	.cin(gnd),
	.combout(\sent_esc~0_combout ),
	.cout());
defparam \sent_esc~0 .lut_mask = 16'hBEFF;
defparam \sent_esc~0 .sum_lutc_input = "datac";

dffeas sent_esc(
	.clk(clk),
	.d(\sent_esc~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sent_esc~q ),
	.prn(vcc));
defparam sent_esc.is_wysiwyg = "true";
defparam sent_esc.power_up = "low";

fiftyfivenm_lcell_comb \in_ready~0 (
	.dataa(\sent_esc~q ),
	.datab(out_data_21),
	.datac(out_data_11),
	.datad(out_data_51),
	.cin(gnd),
	.combout(\in_ready~0_combout ),
	.cout());
defparam \in_ready~0 .lut_mask = 16'hBEFF;
defparam \in_ready~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \in_ready~1 (
	.dataa(out_data_71),
	.datab(out_data_61),
	.datac(out_data_41),
	.datad(out_data_31),
	.cin(gnd),
	.combout(\in_ready~1_combout ),
	.cout());
defparam \in_ready~1 .lut_mask = 16'hBFFF;
defparam \in_ready~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \in_ready~3 (
	.dataa(\in_ready~0_combout ),
	.datab(\in_ready~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_ready~3_combout ),
	.cout());
defparam \in_ready~3 .lut_mask = 16'hEEEE;
defparam \in_ready~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \sent_channel_char~0 (
	.dataa(\always0~0_combout ),
	.datab(\sent_channel_char~q ),
	.datac(\out_data[7]~0_combout ),
	.datad(\in_ready~3_combout ),
	.cin(gnd),
	.combout(\sent_channel_char~0_combout ),
	.cout());
defparam \sent_channel_char~0 .lut_mask = 16'hEFFF;
defparam \sent_channel_char~0 .sum_lutc_input = "datac";

dffeas sent_channel_char(
	.clk(clk),
	.d(\sent_channel_char~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~2_combout ),
	.q(\sent_channel_char~q ),
	.prn(vcc));
defparam sent_channel_char.is_wysiwyg = "true";
defparam sent_channel_char.power_up = "low";

fiftyfivenm_lcell_comb \sent_channel~0 (
	.dataa(\sent_channel_char~q ),
	.datab(out_startofpacket),
	.datac(\stored_channel[0]~q ),
	.datad(\sent_channel~q ),
	.cin(gnd),
	.combout(\sent_channel~0_combout ),
	.cout());
defparam \sent_channel~0 .lut_mask = 16'hEFFF;
defparam \sent_channel~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \sent_channel~1 (
	.dataa(\sent_channel~0_combout ),
	.datab(\sent_channel~q ),
	.datac(\out_data[7]~0_combout ),
	.datad(\in_ready~3_combout ),
	.cin(gnd),
	.combout(\sent_channel~1_combout ),
	.cout());
defparam \sent_channel~1 .lut_mask = 16'hEFFF;
defparam \sent_channel~1 .sum_lutc_input = "datac";

dffeas sent_channel(
	.clk(clk),
	.d(\sent_channel~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_ready~2_combout ),
	.q(\sent_channel~q ),
	.prn(vcc));
defparam sent_channel.is_wysiwyg = "true";
defparam sent_channel.power_up = "low";

fiftyfivenm_lcell_comb \stored_channel[0]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sent_channel~q ),
	.datad(\stored_channel[0]~q ),
	.cin(gnd),
	.combout(\stored_channel[0]~0_combout ),
	.cout());
defparam \stored_channel[0]~0 .lut_mask = 16'hFFF0;
defparam \stored_channel[0]~0 .sum_lutc_input = "datac";

dffeas \stored_channel[0] (
	.clk(clk),
	.d(\stored_channel[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\stored_channel[0]~q ),
	.prn(vcc));
defparam \stored_channel[0] .is_wysiwyg = "true";
defparam \stored_channel[0] .power_up = "low";

fiftyfivenm_lcell_comb \always0~0 (
	.dataa(out_startofpacket),
	.datab(gnd),
	.datac(\stored_channel[0]~q ),
	.datad(\sent_channel~q ),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
defparam \always0~0 .lut_mask = 16'hAFFF;
defparam \always0~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \in_ready~4 (
	.dataa(\in_ready~2_combout ),
	.datab(\sent_sop~q ),
	.datac(out_startofpacket),
	.datad(\always0~0_combout ),
	.cin(gnd),
	.combout(\in_ready~4_combout ),
	.cout());
defparam \in_ready~4 .lut_mask = 16'hEFFF;
defparam \in_ready~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \sent_eop~2 (
	.dataa(out_endofpacket),
	.datab(\sent_eop~q ),
	.datac(\in_ready~4_combout ),
	.datad(\in_ready~3_combout ),
	.cin(gnd),
	.combout(\sent_eop~2_combout ),
	.cout());
defparam \sent_eop~2 .lut_mask = 16'hBEFF;
defparam \sent_eop~2 .sum_lutc_input = "datac";

dffeas sent_eop(
	.clk(clk),
	.d(\sent_eop~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sent_eop~q ),
	.prn(vcc));
defparam sent_eop.is_wysiwyg = "true";
defparam sent_eop.power_up = "low";

fiftyfivenm_lcell_comb \always0~2 (
	.dataa(out_endofpacket),
	.datab(gnd),
	.datac(gnd),
	.datad(\sent_eop~q ),
	.cin(gnd),
	.combout(\always0~2_combout ),
	.cout());
defparam \always0~2 .lut_mask = 16'hAAFF;
defparam \always0~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \sent_sop~3 (
	.dataa(out_startofpacket),
	.datab(\sent_sop~q ),
	.datac(\in_ready~2_combout ),
	.datad(\always0~0_combout ),
	.cin(gnd),
	.combout(\sent_sop~3_combout ),
	.cout());
defparam \sent_sop~3 .lut_mask = 16'hFEFF;
defparam \sent_sop~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \sent_sop~2 (
	.dataa(\always0~2_combout ),
	.datab(\in_ready~3_combout ),
	.datac(\sent_sop~q ),
	.datad(\sent_sop~3_combout ),
	.cin(gnd),
	.combout(\sent_sop~2_combout ),
	.cout());
defparam \sent_sop~2 .lut_mask = 16'hBFFB;
defparam \sent_sop~2 .sum_lutc_input = "datac";

dffeas sent_sop(
	.clk(clk),
	.d(\sent_sop~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sent_sop~q ),
	.prn(vcc));
defparam sent_sop.is_wysiwyg = "true";
defparam sent_sop.power_up = "low";

fiftyfivenm_lcell_comb \out_data[7]~0 (
	.dataa(\sent_sop~q ),
	.datab(\sent_eop~q ),
	.datac(out_endofpacket),
	.datad(out_startofpacket),
	.cin(gnd),
	.combout(\out_data[7]~0_combout ),
	.cout());
defparam \out_data[7]~0 .lut_mask = 16'hEFFF;
defparam \out_data[7]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data[7]~1 (
	.dataa(\out_data[7]~0_combout ),
	.datab(\in_ready~0_combout ),
	.datac(\in_ready~1_combout ),
	.datad(\always0~0_combout ),
	.cin(gnd),
	.combout(\out_data[7]~1_combout ),
	.cout());
defparam \out_data[7]~1 .lut_mask = 16'hFEFF;
defparam \out_data[7]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \always0~1 (
	.dataa(out_startofpacket),
	.datab(gnd),
	.datac(gnd),
	.datad(\sent_sop~q ),
	.cin(gnd),
	.combout(\always0~1_combout ),
	.cout());
defparam \always0~1 .lut_mask = 16'hAAFF;
defparam \always0~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data~2 (
	.dataa(out_data_01),
	.datab(\out_data[7]~1_combout ),
	.datac(\always0~1_combout ),
	.datad(\always0~0_combout ),
	.cin(gnd),
	.combout(\out_data~2_combout ),
	.cout());
defparam \out_data~2 .lut_mask = 16'h8BFF;
defparam \out_data~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_valid~0 (
	.dataa(out_valid2),
	.datab(out_valid1),
	.datac(in_data_toggle),
	.datad(dreg_6),
	.cin(gnd),
	.combout(\out_valid~0_combout ),
	.cout());
defparam \out_valid~0 .lut_mask = 16'hEFFE;
defparam \out_valid~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data~3 (
	.dataa(\out_data[7]~0_combout ),
	.datab(out_data_21),
	.datac(\in_ready~3_combout ),
	.datad(\always0~0_combout ),
	.cin(gnd),
	.combout(\out_data~3_combout ),
	.cout());
defparam \out_data~3 .lut_mask = 16'hEFFF;
defparam \out_data~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data~4 (
	.dataa(\out_data~3_combout ),
	.datab(\always0~0_combout ),
	.datac(gnd),
	.datad(\sent_channel_char~q ),
	.cin(gnd),
	.combout(\out_data~4_combout ),
	.cout());
defparam \out_data~4 .lut_mask = 16'hEEFF;
defparam \out_data~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data~5 (
	.dataa(out_data_11),
	.datab(\out_data[7]~1_combout ),
	.datac(\out_data[7]~0_combout ),
	.datad(\always0~0_combout ),
	.cin(gnd),
	.combout(\out_data~5_combout ),
	.cout());
defparam \out_data~5 .lut_mask = 16'h8BFF;
defparam \out_data~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data~6 (
	.dataa(out_data_61),
	.datab(gnd),
	.datac(\out_data[7]~1_combout ),
	.datad(\sent_channel~0_combout ),
	.cin(gnd),
	.combout(\out_data~6_combout ),
	.cout());
defparam \out_data~6 .lut_mask = 16'hAFFF;
defparam \out_data~6 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data~7 (
	.dataa(out_data_71),
	.datab(\out_data[7]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_data~7_combout ),
	.cout());
defparam \out_data~7 .lut_mask = 16'hEEEE;
defparam \out_data~7 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\sent_esc~q ),
	.datad(out_data_51),
	.cin(gnd),
	.combout(\out_data~8_combout ),
	.cout());
defparam \out_data~8 .lut_mask = 16'h0FF0;
defparam \out_data~8 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data~9 (
	.dataa(\out_data~8_combout ),
	.datab(\out_data[7]~0_combout ),
	.datac(\always0~0_combout ),
	.datad(\sent_channel_char~q ),
	.cin(gnd),
	.combout(\out_data~9_combout ),
	.cout());
defparam \out_data~9 .lut_mask = 16'hA3FF;
defparam \out_data~9 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data~10 (
	.dataa(out_data_31),
	.datab(gnd),
	.datac(\out_data[7]~1_combout ),
	.datad(\sent_channel~0_combout ),
	.cin(gnd),
	.combout(\out_data~10_combout ),
	.cout());
defparam \out_data~10 .lut_mask = 16'hAFFF;
defparam \out_data~10 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \out_data~11 (
	.dataa(out_data_41),
	.datab(gnd),
	.datac(\out_data[7]~1_combout ),
	.datad(\sent_channel~0_combout ),
	.cin(gnd),
	.combout(\out_data~11_combout ),
	.cout());
defparam \out_data~11 .lut_mask = 16'hAFFF;
defparam \out_data~11 .sum_lutc_input = "datac";

endmodule

module ADC_altera_reset_controller (
	altera_reset_synchronizer_int_chain_out,
	clk_clk,
	reset_reset_n)/* synthesis synthesis_greybox=1 */;
output 	altera_reset_synchronizer_int_chain_out;
input 	clk_clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ADC_altera_reset_synchronizer_1 alt_rst_sync_uq1(
	.altera_reset_synchronizer_int_chain_out1(altera_reset_synchronizer_int_chain_out),
	.clk(clk_clk),
	.reset_reset_n(reset_reset_n));

endmodule

module ADC_altera_reset_synchronizer_1 (
	altera_reset_synchronizer_int_chain_out1,
	clk,
	reset_reset_n)/* synthesis synthesis_greybox=1 */;
output 	altera_reset_synchronizer_int_chain_out1;
input 	clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module ADC_ADC_mm_interconnect_0 (
	readdata_0,
	readdata_01,
	read_latency_shift_reg_1,
	src_data_0,
	mem_used_1,
	mem_used_2,
	address_7,
	address_6,
	address_5,
	address_4,
	Equal0,
	address_9,
	address_3,
	address_8,
	hold_waitrequest,
	write,
	av_waitrequest,
	readdata_2,
	readdata_21,
	src_data_2,
	readdata_1,
	readdata_11,
	src_data_1,
	readdata_5,
	src_payload,
	readdata_6,
	src_payload1,
	readdata_4,
	src_payload2,
	readdata_3,
	readdata_31,
	src_data_3,
	readdata_8,
	src_payload3,
	altera_reset_synchronizer_int_chain_out,
	read,
	src1_valid,
	WideOr1,
	write1,
	readdata_10,
	src_payload4,
	readdata_9,
	src_payload5,
	readdata_13,
	src_payload6,
	readdata_15,
	src_payload7,
	readdata_14,
	src_payload8,
	readdata_12,
	src_payload9,
	readdata_111,
	src_payload10,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	readdata_0;
input 	readdata_01;
output 	read_latency_shift_reg_1;
output 	src_data_0;
output 	mem_used_1;
output 	mem_used_2;
input 	address_7;
input 	address_6;
input 	address_5;
input 	address_4;
output 	Equal0;
input 	address_9;
input 	address_3;
input 	address_8;
output 	hold_waitrequest;
input 	write;
output 	av_waitrequest;
input 	readdata_2;
input 	readdata_21;
output 	src_data_2;
input 	readdata_1;
input 	readdata_11;
output 	src_data_1;
input 	readdata_5;
output 	src_payload;
input 	readdata_6;
output 	src_payload1;
input 	readdata_4;
output 	src_payload2;
input 	readdata_3;
input 	readdata_31;
output 	src_data_3;
input 	readdata_8;
output 	src_payload3;
input 	altera_reset_synchronizer_int_chain_out;
input 	read;
output 	src1_valid;
output 	WideOr1;
output 	write1;
input 	readdata_10;
output 	src_payload4;
input 	readdata_9;
output 	src_payload5;
input 	readdata_13;
output 	src_payload6;
input 	readdata_15;
output 	src_payload7;
input 	readdata_14;
output 	src_payload8;
input 	readdata_12;
output 	src_payload9;
input 	readdata_111;
output 	src_payload10;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \adc_sequencer_csr_translator|read_latency_shift_reg[0]~q ;
wire \router|Equal0~1_combout ;
wire \avalonbridge_master_limiter|last_dest_id[0]~q ;
wire \avalonbridge_master_limiter|has_pending_responses~q ;
wire \avalonbridge_master_limiter|suppress_change_dest_id~0_combout ;
wire \avalonbridge_master_agent|av_waitrequest~0_combout ;
wire \adc_sequencer_csr_translator|read_latency_shift_reg~0_combout ;
wire \avalonbridge_master_limiter|last_channel[0]~q ;
wire \adc_sequencer_csr_agent_rsp_fifo|mem[0][103]~q ;
wire \adc_sample_store_csr_agent_rsp_fifo|mem[0][103]~q ;


ADC_altera_avalon_sc_fifo_2 adc_sequencer_csr_agent_rsp_fifo(
	.read_latency_shift_reg_0(\adc_sequencer_csr_translator|read_latency_shift_reg[0]~q ),
	.mem_used_1(mem_used_1),
	.reset(altera_reset_synchronizer_int_chain_out),
	.read(read),
	.src1_valid(src1_valid),
	.read_latency_shift_reg(\adc_sequencer_csr_translator|read_latency_shift_reg~0_combout ),
	.mem_103_0(\adc_sequencer_csr_agent_rsp_fifo|mem[0][103]~q ),
	.clk(clk_clk));

ADC_altera_avalon_sc_fifo_1 adc_sample_store_csr_agent_rsp_fifo(
	.read_latency_shift_reg_1(read_latency_shift_reg_1),
	.mem_used_2(mem_used_2),
	.Equal0(\router|Equal0~1_combout ),
	.hold_waitrequest(hold_waitrequest),
	.has_pending_responses(\avalonbridge_master_limiter|has_pending_responses~q ),
	.write(write),
	.reset(altera_reset_synchronizer_int_chain_out),
	.read(read),
	.last_channel_0(\avalonbridge_master_limiter|last_channel[0]~q ),
	.write1(write1),
	.mem_103_0(\adc_sample_store_csr_agent_rsp_fifo|mem[0][103]~q ),
	.clk(clk_clk));

ADC_altera_merlin_master_agent avalonbridge_master_agent(
	.mem_used_1(mem_used_1),
	.mem_used_2(mem_used_2),
	.Equal0(\router|Equal0~1_combout ),
	.hold_waitrequest1(hold_waitrequest),
	.last_dest_id_0(\avalonbridge_master_limiter|last_dest_id[0]~q ),
	.suppress_change_dest_id(\avalonbridge_master_limiter|suppress_change_dest_id~0_combout ),
	.av_waitrequest(\avalonbridge_master_agent|av_waitrequest~0_combout ),
	.av_waitrequest1(av_waitrequest),
	.altera_reset_synchronizer_int_chain_out(altera_reset_synchronizer_int_chain_out),
	.clk(clk_clk));

ADC_altera_merlin_slave_translator_1 adc_sequencer_csr_translator(
	.read_latency_shift_reg_0(\adc_sequencer_csr_translator|read_latency_shift_reg[0]~q ),
	.mem_used_1(mem_used_1),
	.reset(altera_reset_synchronizer_int_chain_out),
	.read(read),
	.src1_valid(src1_valid),
	.read_latency_shift_reg(\adc_sequencer_csr_translator|read_latency_shift_reg~0_combout ),
	.clk(clk_clk));

ADC_altera_merlin_slave_translator adc_sample_store_csr_translator(
	.read_latency_shift_reg_1(read_latency_shift_reg_1),
	.reset(altera_reset_synchronizer_int_chain_out),
	.write(write1),
	.clk(clk_clk));

ADC_ADC_mm_interconnect_0_rsp_mux rsp_mux(
	.readdata_0(readdata_0),
	.readdata_01(readdata_01),
	.read_latency_shift_reg_0(\adc_sequencer_csr_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_1(read_latency_shift_reg_1),
	.src_data_0(src_data_0),
	.readdata_2(readdata_2),
	.readdata_21(readdata_21),
	.src_data_2(src_data_2),
	.readdata_1(readdata_1),
	.readdata_11(readdata_11),
	.src_data_1(src_data_1),
	.readdata_5(readdata_5),
	.src_payload(src_payload),
	.readdata_6(readdata_6),
	.src_payload1(src_payload1),
	.readdata_4(readdata_4),
	.src_payload2(src_payload2),
	.readdata_3(readdata_3),
	.readdata_31(readdata_31),
	.src_data_3(src_data_3),
	.readdata_8(readdata_8),
	.src_payload3(src_payload3),
	.WideOr11(WideOr1),
	.readdata_10(readdata_10),
	.src_payload4(src_payload4),
	.readdata_9(readdata_9),
	.src_payload5(src_payload5),
	.readdata_13(readdata_13),
	.src_payload6(src_payload6),
	.readdata_15(readdata_15),
	.src_payload7(src_payload7),
	.readdata_14(readdata_14),
	.src_payload8(src_payload8),
	.readdata_12(readdata_12),
	.src_payload9(src_payload9),
	.readdata_111(readdata_111),
	.src_payload10(src_payload10));

ADC_ADC_mm_interconnect_0_cmd_demux cmd_demux(
	.Equal0(\router|Equal0~1_combout ),
	.hold_waitrequest(hold_waitrequest),
	.last_dest_id_0(\avalonbridge_master_limiter|last_dest_id[0]~q ),
	.suppress_change_dest_id(\avalonbridge_master_limiter|suppress_change_dest_id~0_combout ),
	.src1_valid(src1_valid));

ADC_altera_merlin_traffic_limiter avalonbridge_master_limiter(
	.read_latency_shift_reg_0(\adc_sequencer_csr_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg_1(read_latency_shift_reg_1),
	.mem_used_1(mem_used_1),
	.mem_used_2(mem_used_2),
	.cmd_sink_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\router|Equal0~1_combout ,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.last_dest_id_0(\avalonbridge_master_limiter|last_dest_id[0]~q ),
	.has_pending_responses1(\avalonbridge_master_limiter|has_pending_responses~q ),
	.write(write),
	.suppress_change_dest_id(\avalonbridge_master_limiter|suppress_change_dest_id~0_combout ),
	.av_waitrequest(\avalonbridge_master_agent|av_waitrequest~0_combout ),
	.reset(altera_reset_synchronizer_int_chain_out),
	.read(read),
	.last_channel_0(\avalonbridge_master_limiter|last_channel[0]~q ),
	.mem_103_0(\adc_sequencer_csr_agent_rsp_fifo|mem[0][103]~q ),
	.mem_103_01(\adc_sample_store_csr_agent_rsp_fifo|mem[0][103]~q ),
	.clk(clk_clk));

ADC_ADC_mm_interconnect_0_router router(
	.address_7(address_7),
	.address_6(address_6),
	.address_5(address_5),
	.address_4(address_4),
	.Equal0(Equal0),
	.address_9(address_9),
	.address_3(address_3),
	.address_8(address_8),
	.Equal01(\router|Equal0~1_combout ));

endmodule

module ADC_ADC_mm_interconnect_0_cmd_demux (
	Equal0,
	hold_waitrequest,
	last_dest_id_0,
	suppress_change_dest_id,
	src1_valid)/* synthesis synthesis_greybox=1 */;
input 	Equal0;
input 	hold_waitrequest;
input 	last_dest_id_0;
input 	suppress_change_dest_id;
output 	src1_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fiftyfivenm_lcell_comb \src1_valid~0 (
	.dataa(Equal0),
	.datab(hold_waitrequest),
	.datac(last_dest_id_0),
	.datad(suppress_change_dest_id),
	.cin(gnd),
	.combout(src1_valid),
	.cout());
defparam \src1_valid~0 .lut_mask = 16'hFEFF;
defparam \src1_valid~0 .sum_lutc_input = "datac";

endmodule

module ADC_ADC_mm_interconnect_0_router (
	address_7,
	address_6,
	address_5,
	address_4,
	Equal0,
	address_9,
	address_3,
	address_8,
	Equal01)/* synthesis synthesis_greybox=1 */;
input 	address_7;
input 	address_6;
input 	address_5;
input 	address_4;
output 	Equal0;
input 	address_9;
input 	address_3;
input 	address_8;
output 	Equal01;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fiftyfivenm_lcell_comb \Equal0~0 (
	.dataa(address_7),
	.datab(address_6),
	.datac(address_5),
	.datad(address_4),
	.cin(gnd),
	.combout(Equal0),
	.cout());
defparam \Equal0~0 .lut_mask = 16'h7FFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \Equal0~1 (
	.dataa(Equal0),
	.datab(address_9),
	.datac(address_3),
	.datad(address_8),
	.cin(gnd),
	.combout(Equal01),
	.cout());
defparam \Equal0~1 .lut_mask = 16'hEFFF;
defparam \Equal0~1 .sum_lutc_input = "datac";

endmodule

module ADC_ADC_mm_interconnect_0_rsp_mux (
	readdata_0,
	readdata_01,
	read_latency_shift_reg_0,
	read_latency_shift_reg_1,
	src_data_0,
	readdata_2,
	readdata_21,
	src_data_2,
	readdata_1,
	readdata_11,
	src_data_1,
	readdata_5,
	src_payload,
	readdata_6,
	src_payload1,
	readdata_4,
	src_payload2,
	readdata_3,
	readdata_31,
	src_data_3,
	readdata_8,
	src_payload3,
	WideOr11,
	readdata_10,
	src_payload4,
	readdata_9,
	src_payload5,
	readdata_13,
	src_payload6,
	readdata_15,
	src_payload7,
	readdata_14,
	src_payload8,
	readdata_12,
	src_payload9,
	readdata_111,
	src_payload10)/* synthesis synthesis_greybox=1 */;
input 	readdata_0;
input 	readdata_01;
input 	read_latency_shift_reg_0;
input 	read_latency_shift_reg_1;
output 	src_data_0;
input 	readdata_2;
input 	readdata_21;
output 	src_data_2;
input 	readdata_1;
input 	readdata_11;
output 	src_data_1;
input 	readdata_5;
output 	src_payload;
input 	readdata_6;
output 	src_payload1;
input 	readdata_4;
output 	src_payload2;
input 	readdata_3;
input 	readdata_31;
output 	src_data_3;
input 	readdata_8;
output 	src_payload3;
output 	WideOr11;
input 	readdata_10;
output 	src_payload4;
input 	readdata_9;
output 	src_payload5;
input 	readdata_13;
output 	src_payload6;
input 	readdata_15;
output 	src_payload7;
input 	readdata_14;
output 	src_payload8;
input 	readdata_12;
output 	src_payload9;
input 	readdata_111;
output 	src_payload10;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



fiftyfivenm_lcell_comb \src_data[0] (
	.dataa(readdata_0),
	.datab(readdata_01),
	.datac(read_latency_shift_reg_0),
	.datad(read_latency_shift_reg_1),
	.cin(gnd),
	.combout(src_data_0),
	.cout());
defparam \src_data[0] .lut_mask = 16'hFFFE;
defparam \src_data[0] .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \src_data[2] (
	.dataa(read_latency_shift_reg_1),
	.datab(read_latency_shift_reg_0),
	.datac(readdata_2),
	.datad(readdata_21),
	.cin(gnd),
	.combout(src_data_2),
	.cout());
defparam \src_data[2] .lut_mask = 16'hFFFE;
defparam \src_data[2] .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \src_data[1] (
	.dataa(read_latency_shift_reg_1),
	.datab(read_latency_shift_reg_0),
	.datac(readdata_1),
	.datad(readdata_11),
	.cin(gnd),
	.combout(src_data_1),
	.cout());
defparam \src_data[1] .lut_mask = 16'hFFFE;
defparam \src_data[1] .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \src_payload~0 (
	.dataa(read_latency_shift_reg_1),
	.datab(readdata_5),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload),
	.cout());
defparam \src_payload~0 .lut_mask = 16'hEEEE;
defparam \src_payload~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \src_payload~1 (
	.dataa(read_latency_shift_reg_1),
	.datab(readdata_6),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload1),
	.cout());
defparam \src_payload~1 .lut_mask = 16'hEEEE;
defparam \src_payload~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \src_payload~2 (
	.dataa(read_latency_shift_reg_1),
	.datab(readdata_4),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload2),
	.cout());
defparam \src_payload~2 .lut_mask = 16'hEEEE;
defparam \src_payload~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \src_data[3] (
	.dataa(read_latency_shift_reg_1),
	.datab(read_latency_shift_reg_0),
	.datac(readdata_3),
	.datad(readdata_31),
	.cin(gnd),
	.combout(src_data_3),
	.cout());
defparam \src_data[3] .lut_mask = 16'hFFFE;
defparam \src_data[3] .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \src_payload~3 (
	.dataa(read_latency_shift_reg_1),
	.datab(readdata_8),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload3),
	.cout());
defparam \src_payload~3 .lut_mask = 16'hEEEE;
defparam \src_payload~3 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb WideOr1(
	.dataa(read_latency_shift_reg_1),
	.datab(read_latency_shift_reg_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(WideOr11),
	.cout());
defparam WideOr1.lut_mask = 16'hEEEE;
defparam WideOr1.sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \src_payload~4 (
	.dataa(read_latency_shift_reg_1),
	.datab(readdata_10),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload4),
	.cout());
defparam \src_payload~4 .lut_mask = 16'hEEEE;
defparam \src_payload~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \src_payload~5 (
	.dataa(read_latency_shift_reg_1),
	.datab(readdata_9),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload5),
	.cout());
defparam \src_payload~5 .lut_mask = 16'hEEEE;
defparam \src_payload~5 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \src_payload~6 (
	.dataa(read_latency_shift_reg_1),
	.datab(readdata_13),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload6),
	.cout());
defparam \src_payload~6 .lut_mask = 16'hEEEE;
defparam \src_payload~6 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \src_payload~7 (
	.dataa(read_latency_shift_reg_1),
	.datab(readdata_15),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload7),
	.cout());
defparam \src_payload~7 .lut_mask = 16'hEEEE;
defparam \src_payload~7 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \src_payload~8 (
	.dataa(read_latency_shift_reg_1),
	.datab(readdata_14),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload8),
	.cout());
defparam \src_payload~8 .lut_mask = 16'hEEEE;
defparam \src_payload~8 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \src_payload~9 (
	.dataa(read_latency_shift_reg_1),
	.datab(readdata_12),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload9),
	.cout());
defparam \src_payload~9 .lut_mask = 16'hEEEE;
defparam \src_payload~9 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \src_payload~10 (
	.dataa(read_latency_shift_reg_1),
	.datab(readdata_111),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(src_payload10),
	.cout());
defparam \src_payload~10 .lut_mask = 16'hEEEE;
defparam \src_payload~10 .sum_lutc_input = "datac";

endmodule

module ADC_altera_avalon_sc_fifo_1 (
	read_latency_shift_reg_1,
	mem_used_2,
	Equal0,
	hold_waitrequest,
	has_pending_responses,
	write,
	reset,
	read,
	last_channel_0,
	write1,
	mem_103_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	read_latency_shift_reg_1;
output 	mem_used_2;
input 	Equal0;
input 	hold_waitrequest;
input 	has_pending_responses;
input 	write;
input 	reset;
input 	read;
input 	last_channel_0;
output 	write1;
output 	mem_103_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~4_combout ;
wire \mem_used[0]~5_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~3_combout ;
wire \mem_used[1]~q ;
wire \read~0_combout ;
wire \mem_used[2]~2_combout ;
wire \write~0_combout ;
wire \mem[2][103]~q ;
wire \mem~2_combout ;
wire \mem[1][103]~3_combout ;
wire \mem[1][103]~q ;
wire \mem[0][103]~0_combout ;
wire \mem[0][103]~1_combout ;


dffeas \mem_used[2] (
	.clk(clk),
	.d(\mem_used[2]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_2),
	.prn(vcc));
defparam \mem_used[2] .is_wysiwyg = "true";
defparam \mem_used[2] .power_up = "low";

fiftyfivenm_lcell_comb \write~1 (
	.dataa(hold_waitrequest),
	.datab(\write~0_combout ),
	.datac(Equal0),
	.datad(mem_used_2),
	.cin(gnd),
	.combout(write1),
	.cout());
defparam \write~1 .lut_mask = 16'hEFFF;
defparam \write~1 .sum_lutc_input = "datac";

dffeas \mem[0][103] (
	.clk(clk),
	.d(\mem[0][103]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_103_0),
	.prn(vcc));
defparam \mem[0][103] .is_wysiwyg = "true";
defparam \mem[0][103] .power_up = "low";

fiftyfivenm_lcell_comb \mem_used[0]~4 (
	.dataa(write1),
	.datab(\mem_used[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_used[0]~4_combout ),
	.cout());
defparam \mem_used[0]~4 .lut_mask = 16'hEEEE;
defparam \mem_used[0]~4 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \mem_used[0]~5 (
	.dataa(read_latency_shift_reg_1),
	.datab(\mem_used[0]~q ),
	.datac(write1),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_used[0]~5_combout ),
	.cout());
defparam \mem_used[0]~5 .lut_mask = 16'h9696;
defparam \mem_used[0]~5 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[0]~5_combout ),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

fiftyfivenm_lcell_comb \mem_used[1]~3 (
	.dataa(mem_used_2),
	.datab(\mem_used[0]~q ),
	.datac(write1),
	.datad(gnd),
	.cin(gnd),
	.combout(\mem_used[1]~3_combout ),
	.cout());
defparam \mem_used[1]~3 .lut_mask = 16'hFEFE;
defparam \mem_used[1]~3 .sum_lutc_input = "datac";

dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[0]~5_combout ),
	.q(\mem_used[1]~q ),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

fiftyfivenm_lcell_comb \read~0 (
	.dataa(read_latency_shift_reg_1),
	.datab(\mem_used[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\read~0_combout ),
	.cout());
defparam \read~0 .lut_mask = 16'hEEEE;
defparam \read~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \mem_used[2]~2 (
	.dataa(mem_used_2),
	.datab(write1),
	.datac(\mem_used[1]~q ),
	.datad(\read~0_combout ),
	.cin(gnd),
	.combout(\mem_used[2]~2_combout ),
	.cout());
defparam \mem_used[2]~2 .lut_mask = 16'hFBFE;
defparam \mem_used[2]~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \write~0 (
	.dataa(read),
	.datab(write),
	.datac(last_channel_0),
	.datad(has_pending_responses),
	.cin(gnd),
	.combout(\write~0_combout ),
	.cout());
defparam \write~0 .lut_mask = 16'hFEFF;
defparam \write~0 .sum_lutc_input = "datac";

dffeas \mem[2][103] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[2][103]~q ),
	.prn(vcc));
defparam \mem[2][103] .is_wysiwyg = "true";
defparam \mem[2][103] .power_up = "low";

fiftyfivenm_lcell_comb \mem~2 (
	.dataa(\mem[2][103]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(mem_used_2),
	.cin(gnd),
	.combout(\mem~2_combout ),
	.cout());
defparam \mem~2 .lut_mask = 16'hAAFF;
defparam \mem~2 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \mem[1][103]~3 (
	.dataa(\mem~2_combout ),
	.datab(\mem[1][103]~q ),
	.datac(\mem_used[1]~q ),
	.datad(\read~0_combout ),
	.cin(gnd),
	.combout(\mem[1][103]~3_combout ),
	.cout());
defparam \mem[1][103]~3 .lut_mask = 16'hEFFE;
defparam \mem[1][103]~3 .sum_lutc_input = "datac";

dffeas \mem[1][103] (
	.clk(clk),
	.d(\mem[1][103]~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][103]~q ),
	.prn(vcc));
defparam \mem[1][103] .is_wysiwyg = "true";
defparam \mem[1][103] .power_up = "low";

fiftyfivenm_lcell_comb \mem[0][103]~0 (
	.dataa(\mem_used[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(read_latency_shift_reg_1),
	.cin(gnd),
	.combout(\mem[0][103]~0_combout ),
	.cout());
defparam \mem[0][103]~0 .lut_mask = 16'hAAFF;
defparam \mem[0][103]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \mem[0][103]~1 (
	.dataa(mem_103_0),
	.datab(\mem[1][103]~q ),
	.datac(\mem_used[1]~q ),
	.datad(\mem[0][103]~0_combout ),
	.cin(gnd),
	.combout(\mem[0][103]~1_combout ),
	.cout());
defparam \mem[0][103]~1 .lut_mask = 16'hAFCF;
defparam \mem[0][103]~1 .sum_lutc_input = "datac";

endmodule

module ADC_altera_avalon_sc_fifo_2 (
	read_latency_shift_reg_0,
	mem_used_1,
	reset,
	read,
	src1_valid,
	read_latency_shift_reg,
	mem_103_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	read_latency_shift_reg_0;
output 	mem_used_1;
input 	reset;
input 	read;
input 	src1_valid;
input 	read_latency_shift_reg;
output 	mem_103_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~2_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem[1][103]~q ;
wire \mem~0_combout ;
wire \mem[0][103]~1_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][103] (
	.clk(clk),
	.d(\mem[0][103]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_103_0),
	.prn(vcc));
defparam \mem[0][103] .is_wysiwyg = "true";
defparam \mem[0][103] .power_up = "low";

fiftyfivenm_lcell_comb \mem_used[0]~2 (
	.dataa(read_latency_shift_reg),
	.datab(\mem_used[0]~q ),
	.datac(mem_used_1),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[0]~2_combout ),
	.cout());
defparam \mem_used[0]~2 .lut_mask = 16'hFEFF;
defparam \mem_used[0]~2 .sum_lutc_input = "datac";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

fiftyfivenm_lcell_comb \mem_used[1]~0 (
	.dataa(read),
	.datab(src1_valid),
	.datac(\mem_used[0]~q ),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem_used[1]~0_combout ),
	.cout());
defparam \mem_used[1]~0 .lut_mask = 16'hFEFF;
defparam \mem_used[1]~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \mem_used[1]~1 (
	.dataa(\mem_used[1]~0_combout ),
	.datab(mem_used_1),
	.datac(read_latency_shift_reg_0),
	.datad(\mem_used[0]~q ),
	.cin(gnd),
	.combout(\mem_used[1]~1_combout ),
	.cout());
defparam \mem_used[1]~1 .lut_mask = 16'hEFFF;
defparam \mem_used[1]~1 .sum_lutc_input = "datac";

dffeas \mem[1][103] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][103]~q ),
	.prn(vcc));
defparam \mem[1][103] .is_wysiwyg = "true";
defparam \mem[1][103] .power_up = "low";

fiftyfivenm_lcell_comb \mem~0 (
	.dataa(\mem[1][103]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\mem~0_combout ),
	.cout());
defparam \mem~0 .lut_mask = 16'hAAFF;
defparam \mem~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \mem[0][103]~1 (
	.dataa(\mem~0_combout ),
	.datab(mem_103_0),
	.datac(\mem_used[0]~q ),
	.datad(read_latency_shift_reg_0),
	.cin(gnd),
	.combout(\mem[0][103]~1_combout ),
	.cout());
defparam \mem[0][103]~1 .lut_mask = 16'hEFFE;
defparam \mem[0][103]~1 .sum_lutc_input = "datac";

endmodule

module ADC_altera_merlin_master_agent (
	mem_used_1,
	mem_used_2,
	Equal0,
	hold_waitrequest1,
	last_dest_id_0,
	suppress_change_dest_id,
	av_waitrequest,
	av_waitrequest1,
	altera_reset_synchronizer_int_chain_out,
	clk)/* synthesis synthesis_greybox=1 */;
input 	mem_used_1;
input 	mem_used_2;
input 	Equal0;
output 	hold_waitrequest1;
input 	last_dest_id_0;
input 	suppress_change_dest_id;
output 	av_waitrequest;
output 	av_waitrequest1;
input 	altera_reset_synchronizer_int_chain_out;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas hold_waitrequest(
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(altera_reset_synchronizer_int_chain_out),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(hold_waitrequest1),
	.prn(vcc));
defparam hold_waitrequest.is_wysiwyg = "true";
defparam hold_waitrequest.power_up = "low";

fiftyfivenm_lcell_comb \av_waitrequest~0 (
	.dataa(hold_waitrequest1),
	.datab(Equal0),
	.datac(last_dest_id_0),
	.datad(suppress_change_dest_id),
	.cin(gnd),
	.combout(av_waitrequest),
	.cout());
defparam \av_waitrequest~0 .lut_mask = 16'hBEFF;
defparam \av_waitrequest~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \av_waitrequest~1 (
	.dataa(mem_used_1),
	.datab(mem_used_2),
	.datac(Equal0),
	.datad(av_waitrequest),
	.cin(gnd),
	.combout(av_waitrequest1),
	.cout());
defparam \av_waitrequest~1 .lut_mask = 16'hACFF;
defparam \av_waitrequest~1 .sum_lutc_input = "datac";

endmodule

module ADC_altera_merlin_slave_translator (
	read_latency_shift_reg_1,
	reset,
	write,
	clk)/* synthesis synthesis_greybox=1 */;
output 	read_latency_shift_reg_1;
input 	reset;
input 	write;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg[0]~q ;


dffeas \read_latency_shift_reg[1] (
	.clk(clk),
	.d(\read_latency_shift_reg[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_1),
	.prn(vcc));
defparam \read_latency_shift_reg[1] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[1] .power_up = "low";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(write),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read_latency_shift_reg[0]~q ),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

endmodule

module ADC_altera_merlin_slave_translator_1 (
	read_latency_shift_reg_0,
	mem_used_1,
	reset,
	read,
	src1_valid,
	read_latency_shift_reg,
	clk)/* synthesis synthesis_greybox=1 */;
output 	read_latency_shift_reg_0;
input 	mem_used_1;
input 	reset;
input 	read;
input 	src1_valid;
output 	read_latency_shift_reg;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(read_latency_shift_reg),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

fiftyfivenm_lcell_comb \read_latency_shift_reg~0 (
	.dataa(read),
	.datab(src1_valid),
	.datac(gnd),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(read_latency_shift_reg),
	.cout());
defparam \read_latency_shift_reg~0 .lut_mask = 16'hEEFF;
defparam \read_latency_shift_reg~0 .sum_lutc_input = "datac";

endmodule

module ADC_altera_merlin_traffic_limiter (
	read_latency_shift_reg_0,
	read_latency_shift_reg_1,
	mem_used_1,
	mem_used_2,
	cmd_sink_data,
	last_dest_id_0,
	has_pending_responses1,
	write,
	suppress_change_dest_id,
	av_waitrequest,
	reset,
	read,
	last_channel_0,
	mem_103_0,
	mem_103_01,
	clk)/* synthesis synthesis_greybox=1 */;
input 	read_latency_shift_reg_0;
input 	read_latency_shift_reg_1;
input 	mem_used_1;
input 	mem_used_2;
input 	[101:0] cmd_sink_data;
output 	last_dest_id_0;
output 	has_pending_responses1;
input 	write;
output 	suppress_change_dest_id;
input 	av_waitrequest;
input 	reset;
input 	read;
output 	last_channel_0;
input 	mem_103_0;
input 	mem_103_01;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \save_dest_id~0_combout ;
wire \response_sink_accepted~0_combout ;
wire \nonposted_cmd_accepted~0_combout ;
wire \pending_response_count[0]~1_combout ;
wire \pending_response_count[1]~0_combout ;
wire \pending_response_count[0]~q ;
wire \Add0~0_combout ;
wire \pending_response_count[1]~q ;
wire \has_pending_responses~0_combout ;
wire \has_pending_responses~1_combout ;
wire \last_channel[0]~0_combout ;


dffeas \last_dest_id[0] (
	.clk(clk),
	.d(cmd_sink_data[88]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_dest_id_0),
	.prn(vcc));
defparam \last_dest_id[0] .is_wysiwyg = "true";
defparam \last_dest_id[0] .power_up = "low";

dffeas has_pending_responses(
	.clk(clk),
	.d(\has_pending_responses~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(has_pending_responses1),
	.prn(vcc));
defparam has_pending_responses.is_wysiwyg = "true";
defparam has_pending_responses.power_up = "low";

fiftyfivenm_lcell_comb \suppress_change_dest_id~0 (
	.dataa(has_pending_responses1),
	.datab(gnd),
	.datac(gnd),
	.datad(write),
	.cin(gnd),
	.combout(suppress_change_dest_id),
	.cout());
defparam \suppress_change_dest_id~0 .lut_mask = 16'hAAFF;
defparam \suppress_change_dest_id~0 .sum_lutc_input = "datac";

dffeas \last_channel[0] (
	.clk(clk),
	.d(\last_channel[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_channel_0),
	.prn(vcc));
defparam \last_channel[0] .is_wysiwyg = "true";
defparam \last_channel[0] .power_up = "low";

fiftyfivenm_lcell_comb \save_dest_id~0 (
	.dataa(av_waitrequest),
	.datab(read),
	.datac(gnd),
	.datad(write),
	.cin(gnd),
	.combout(\save_dest_id~0_combout ),
	.cout());
defparam \save_dest_id~0 .lut_mask = 16'hEEFF;
defparam \save_dest_id~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \response_sink_accepted~0 (
	.dataa(read_latency_shift_reg_1),
	.datab(read_latency_shift_reg_0),
	.datac(mem_103_0),
	.datad(mem_103_01),
	.cin(gnd),
	.combout(\response_sink_accepted~0_combout ),
	.cout());
defparam \response_sink_accepted~0 .lut_mask = 16'hFFFE;
defparam \response_sink_accepted~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \nonposted_cmd_accepted~0 (
	.dataa(\save_dest_id~0_combout ),
	.datab(cmd_sink_data[88]),
	.datac(mem_used_2),
	.datad(mem_used_1),
	.cin(gnd),
	.combout(\nonposted_cmd_accepted~0_combout ),
	.cout());
defparam \nonposted_cmd_accepted~0 .lut_mask = 16'h8BFF;
defparam \nonposted_cmd_accepted~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \pending_response_count[0]~1 (
	.dataa(\pending_response_count[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\pending_response_count[0]~1_combout ),
	.cout());
defparam \pending_response_count[0]~1 .lut_mask = 16'h5555;
defparam \pending_response_count[0]~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \pending_response_count[1]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\nonposted_cmd_accepted~0_combout ),
	.datad(\response_sink_accepted~0_combout ),
	.cin(gnd),
	.combout(\pending_response_count[1]~0_combout ),
	.cout());
defparam \pending_response_count[1]~0 .lut_mask = 16'h0FF0;
defparam \pending_response_count[1]~0 .sum_lutc_input = "datac";

dffeas \pending_response_count[0] (
	.clk(clk),
	.d(\pending_response_count[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pending_response_count[1]~0_combout ),
	.q(\pending_response_count[0]~q ),
	.prn(vcc));
defparam \pending_response_count[0] .is_wysiwyg = "true";
defparam \pending_response_count[0] .power_up = "low";

fiftyfivenm_lcell_comb \Add0~0 (
	.dataa(\response_sink_accepted~0_combout ),
	.datab(\pending_response_count[1]~q ),
	.datac(\pending_response_count[0]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout());
defparam \Add0~0 .lut_mask = 16'h9696;
defparam \Add0~0 .sum_lutc_input = "datac";

dffeas \pending_response_count[1] (
	.clk(clk),
	.d(\Add0~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\pending_response_count[1]~0_combout ),
	.q(\pending_response_count[1]~q ),
	.prn(vcc));
defparam \pending_response_count[1] .is_wysiwyg = "true";
defparam \pending_response_count[1] .power_up = "low";

fiftyfivenm_lcell_comb \has_pending_responses~0 (
	.dataa(\pending_response_count[1]~q ),
	.datab(\pending_response_count[0]~q ),
	.datac(has_pending_responses1),
	.datad(gnd),
	.cin(gnd),
	.combout(\has_pending_responses~0_combout ),
	.cout());
defparam \has_pending_responses~0 .lut_mask = 16'h8D8D;
defparam \has_pending_responses~0 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \has_pending_responses~1 (
	.dataa(\response_sink_accepted~0_combout ),
	.datab(\nonposted_cmd_accepted~0_combout ),
	.datac(has_pending_responses1),
	.datad(\has_pending_responses~0_combout ),
	.cin(gnd),
	.combout(\has_pending_responses~1_combout ),
	.cout());
defparam \has_pending_responses~1 .lut_mask = 16'hFDFF;
defparam \has_pending_responses~1 .sum_lutc_input = "datac";

fiftyfivenm_lcell_comb \last_channel[0]~0 (
	.dataa(cmd_sink_data[88]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\last_channel[0]~0_combout ),
	.cout());
defparam \last_channel[0]~0 .lut_mask = 16'h5555;
defparam \last_channel[0]~0 .sum_lutc_input = "datac";

endmodule

module ADC_ADC_PLL (
	wire_pll7_locked,
	wire_pll7_clk_0,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	wire_pll7_locked;
output 	wire_pll7_clk_0;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ADC_ADC_PLL_altpll_5q22 sd1(
	.wire_pll7_locked(wire_pll7_locked),
	.clk({clk_unconnected_wire_4,clk_unconnected_wire_3,clk_unconnected_wire_2,clk_unconnected_wire_1,wire_pll7_clk_0}),
	.inclk({gnd,clk_clk}));

endmodule

module ADC_ADC_PLL_altpll_5q22 (
	wire_pll7_locked,
	clk,
	inclk)/* synthesis synthesis_greybox=1 */;
output 	wire_pll7_locked;
output 	[4:0] clk;
input 	[1:0] inclk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wire_pll7_clk[1] ;
wire \wire_pll7_clk[2] ;
wire \wire_pll7_clk[3] ;
wire \wire_pll7_clk[4] ;
wire wire_pll7_fbout;

wire [4:0] pll7_CLK_bus;

assign clk[0] = pll7_CLK_bus[0];
assign \wire_pll7_clk[1]  = pll7_CLK_bus[1];
assign \wire_pll7_clk[2]  = pll7_CLK_bus[2];
assign \wire_pll7_clk[3]  = pll7_CLK_bus[3];
assign \wire_pll7_clk[4]  = pll7_CLK_bus[4];

fiftyfivenm_pll pll7(
	.areset(gnd),
	.pfdena(vcc),
	.fbin(wire_pll7_fbout),
	.phaseupdown(gnd),
	.phasestep(gnd),
	.scandata(gnd),
	.scanclk(gnd),
	.scanclkena(vcc),
	.configupdate(gnd),
	.clkswitch(gnd),
	.inclk({gnd,inclk[0]}),
	.phasecounterselect(3'b000),
	.phasedone(),
	.scandataout(),
	.scandone(),
	.activeclock(),
	.locked(wire_pll7_locked),
	.vcooverrange(),
	.vcounderrange(),
	.fbout(wire_pll7_fbout),
	.clk(pll7_CLK_bus),
	.clkbad());
defparam pll7.auto_settings = "false";
defparam pll7.bandwidth_type = "auto";
defparam pll7.c0_high = 40;
defparam pll7.c0_initial = 1;
defparam pll7.c0_low = 40;
defparam pll7.c0_mode = "even";
defparam pll7.c0_ph = 0;
defparam pll7.c1_high = 1;
defparam pll7.c1_initial = 1;
defparam pll7.c1_low = 1;
defparam pll7.c1_mode = "bypass";
defparam pll7.c1_ph = 0;
defparam pll7.c1_use_casc_in = "off";
defparam pll7.c2_high = 1;
defparam pll7.c2_initial = 1;
defparam pll7.c2_low = 1;
defparam pll7.c2_mode = "bypass";
defparam pll7.c2_ph = 0;
defparam pll7.c2_use_casc_in = "off";
defparam pll7.c3_high = 1;
defparam pll7.c3_initial = 1;
defparam pll7.c3_low = 1;
defparam pll7.c3_mode = "bypass";
defparam pll7.c3_ph = 0;
defparam pll7.c3_use_casc_in = "off";
defparam pll7.c4_high = 1;
defparam pll7.c4_initial = 1;
defparam pll7.c4_low = 1;
defparam pll7.c4_mode = "bypass";
defparam pll7.c4_ph = 0;
defparam pll7.c4_use_casc_in = "off";
defparam pll7.charge_pump_current_bits = 2;
defparam pll7.clk0_counter = "c0";
defparam pll7.clk0_divide_by = 5;
defparam pll7.clk0_duty_cycle = 50;
defparam pll7.clk0_multiply_by = 1;
defparam pll7.clk0_phase_shift = "0";
defparam pll7.clk1_counter = "unused";
defparam pll7.clk1_divide_by = 0;
defparam pll7.clk1_duty_cycle = 50;
defparam pll7.clk1_multiply_by = 0;
defparam pll7.clk1_phase_shift = "0";
defparam pll7.clk2_counter = "unused";
defparam pll7.clk2_divide_by = 0;
defparam pll7.clk2_duty_cycle = 50;
defparam pll7.clk2_multiply_by = 0;
defparam pll7.clk2_phase_shift = "0";
defparam pll7.clk3_counter = "unused";
defparam pll7.clk3_divide_by = 0;
defparam pll7.clk3_duty_cycle = 50;
defparam pll7.clk3_multiply_by = 0;
defparam pll7.clk3_phase_shift = "0";
defparam pll7.clk4_counter = "unused";
defparam pll7.clk4_divide_by = 0;
defparam pll7.clk4_duty_cycle = 50;
defparam pll7.clk4_multiply_by = 0;
defparam pll7.clk4_phase_shift = "0";
defparam pll7.compensate_clock = "clock0";
defparam pll7.inclk0_input_frequency = 20000;
defparam pll7.inclk1_input_frequency = 0;
defparam pll7.loop_filter_c_bits = 2;
defparam pll7.loop_filter_r_bits = 1;
defparam pll7.m = 16;
defparam pll7.m_initial = 1;
defparam pll7.m_ph = 0;
defparam pll7.n = 1;
defparam pll7.operation_mode = "normal";
defparam pll7.pfd_max = 0;
defparam pll7.pfd_min = 0;
defparam pll7.self_reset_on_loss_lock = "off";
defparam pll7.simulation_type = "timing";
defparam pll7.switch_over_type = "auto";
defparam pll7.vco_center = 0;
defparam pll7.vco_divide_by = 0;
defparam pll7.vco_frequency_control = "auto";
defparam pll7.vco_max = 0;
defparam pll7.vco_min = 0;
defparam pll7.vco_multiply_by = 0;
defparam pll7.vco_phase_shift_step = 0;
defparam pll7.vco_post_scale = 1;

endmodule

module ADC_altera_reset_controller_1 (
	altera_reset_synchronizer_int_chain_out,
	clk_clk,
	reset_reset_n)/* synthesis synthesis_greybox=1 */;
output 	altera_reset_synchronizer_int_chain_out;
input 	clk_clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ADC_altera_reset_synchronizer_3 alt_rst_sync_uq1(
	.altera_reset_synchronizer_int_chain_out1(altera_reset_synchronizer_int_chain_out),
	.clk(clk_clk),
	.reset_reset_n(reset_reset_n));

endmodule

module ADC_altera_reset_synchronizer_3 (
	altera_reset_synchronizer_int_chain_out1,
	clk,
	reset_reset_n)/* synthesis synthesis_greybox=1 */;
output 	altera_reset_synchronizer_int_chain_out1;
input 	clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule
